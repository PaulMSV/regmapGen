// Created with regmapGen v1.0.3

Uchip_regmap0 Uchip_regmap0_wrapper(
    // System
    .clk(clk),
    .rst(rst),

    // DisDrvConfig0.DDIS_DRVB_CFG_INJ
    .disdrvconfig0_ddis_drvb_cfg_inj_en(disdrvconfig0_ddis_drvb_cfg_inj_en),
    .disdrvconfig0_ddis_drvb_cfg_inj_in(disdrvconfig0_ddis_drvb_cfg_inj_in),
    .disdrvconfig0_ddis_drvb_cfg_inj_out(disdrvconfig0_ddis_drvb_cfg_inj_out),
    // DisDrvConfig0.DDIS_DRVB_CFG_IGN
    .disdrvconfig0_ddis_drvb_cfg_ign_en(disdrvconfig0_ddis_drvb_cfg_ign_en),
    .disdrvconfig0_ddis_drvb_cfg_ign_in(disdrvconfig0_ddis_drvb_cfg_ign_in),
    .disdrvconfig0_ddis_drvb_cfg_ign_out(disdrvconfig0_ddis_drvb_cfg_ign_out),

    // DisDrvConfig1.DDIS_DRVB_CFG_RLY
    .disdrvconfig1_ddis_drvb_cfg_rly_en(disdrvconfig1_ddis_drvb_cfg_rly_en),
    .disdrvconfig1_ddis_drvb_cfg_rly_in(disdrvconfig1_ddis_drvb_cfg_rly_in),
    .disdrvconfig1_ddis_drvb_cfg_rly_out(disdrvconfig1_ddis_drvb_cfg_rly_out),

    // DisDrvConfig2.DDIS_DRVB_CFG_RLY
    .disdrvconfig2_ddis_drvb_cfg_rly_en(disdrvconfig2_ddis_drvb_cfg_rly_en),
    .disdrvconfig2_ddis_drvb_cfg_rly_in(disdrvconfig2_ddis_drvb_cfg_rly_in),
    .disdrvconfig2_ddis_drvb_cfg_rly_out(disdrvconfig2_ddis_drvb_cfg_rly_out),
    // DisDrvConfig2.DDIS_DRVB_CFG_VLV
    .disdrvconfig2_ddis_drvb_cfg_vlv_en(disdrvconfig2_ddis_drvb_cfg_vlv_en),
    .disdrvconfig2_ddis_drvb_cfg_vlv_in(disdrvconfig2_ddis_drvb_cfg_vlv_in),
    .disdrvconfig2_ddis_drvb_cfg_vlv_out(disdrvconfig2_ddis_drvb_cfg_vlv_out),
    // DisDrvConfig2.DDIS_DRVB_CFG_HTR
    .disdrvconfig2_ddis_drvb_cfg_htr_en(disdrvconfig2_ddis_drvb_cfg_htr_en),
    .disdrvconfig2_ddis_drvb_cfg_htr_in(disdrvconfig2_ddis_drvb_cfg_htr_in),
    .disdrvconfig2_ddis_drvb_cfg_htr_out(disdrvconfig2_ddis_drvb_cfg_htr_out),
    // DisDrvConfig2.DDIS_DRVB_CFG_HB
    .disdrvconfig2_ddis_drvb_cfg_hb_en(disdrvconfig2_ddis_drvb_cfg_hb_en),
    .disdrvconfig2_ddis_drvb_cfg_hb_in(disdrvconfig2_ddis_drvb_cfg_hb_in),
    .disdrvconfig2_ddis_drvb_cfg_hb_out(disdrvconfig2_ddis_drvb_cfg_hb_out),

    // DenConfig0.DEN_DRV_CFG_IGN
    .denconfig0_den_drv_cfg_ign_en(denconfig0_den_drv_cfg_ign_en),
    .denconfig0_den_drv_cfg_ign_in(denconfig0_den_drv_cfg_ign_in),
    .denconfig0_den_drv_cfg_ign_out(denconfig0_den_drv_cfg_ign_out),

    // DenConfig1.DEN_DRV_CFG_RLY1
    .denconfig1_den_drv_cfg_rly1_en(denconfig1_den_drv_cfg_rly1_en),
    .denconfig1_den_drv_cfg_rly1_in(denconfig1_den_drv_cfg_rly1_in),
    .denconfig1_den_drv_cfg_rly1_out(denconfig1_den_drv_cfg_rly1_out),
    // DenConfig1.DEN_RLY_CFG_RLY1
    .denconfig1_den_rly_cfg_rly1_en(denconfig1_den_rly_cfg_rly1_en),
    .denconfig1_den_rly_cfg_rly1_in(denconfig1_den_rly_cfg_rly1_in),
    .denconfig1_den_rly_cfg_rly1_out(denconfig1_den_rly_cfg_rly1_out),
    // DenConfig1.DEN_DRV_CFG_RLY2
    .denconfig1_den_drv_cfg_rly2_en(denconfig1_den_drv_cfg_rly2_en),
    .denconfig1_den_drv_cfg_rly2_in(denconfig1_den_drv_cfg_rly2_in),
    .denconfig1_den_drv_cfg_rly2_out(denconfig1_den_drv_cfg_rly2_out),
    // DenConfig1.DEN_RLY_CFG_RLY2
    .denconfig1_den_rly_cfg_rly2_en(denconfig1_den_rly_cfg_rly2_en),
    .denconfig1_den_rly_cfg_rly2_in(denconfig1_den_rly_cfg_rly2_in),
    .denconfig1_den_rly_cfg_rly2_out(denconfig1_den_rly_cfg_rly2_out),
    // DenConfig1.DEN_DRV_CFG_RLY3
    .denconfig1_den_drv_cfg_rly3_en(denconfig1_den_drv_cfg_rly3_en),
    .denconfig1_den_drv_cfg_rly3_in(denconfig1_den_drv_cfg_rly3_in),
    .denconfig1_den_drv_cfg_rly3_out(denconfig1_den_drv_cfg_rly3_out),
    // DenConfig1.DEN_RLY_CFG_RLY3
    .denconfig1_den_rly_cfg_rly3_en(denconfig1_den_rly_cfg_rly3_en),
    .denconfig1_den_rly_cfg_rly3_in(denconfig1_den_rly_cfg_rly3_in),
    .denconfig1_den_rly_cfg_rly3_out(denconfig1_den_rly_cfg_rly3_out),
    // DenConfig1.DEN_DRV_CFG_RLY4
    .denconfig1_den_drv_cfg_rly4_en(denconfig1_den_drv_cfg_rly4_en),
    .denconfig1_den_drv_cfg_rly4_in(denconfig1_den_drv_cfg_rly4_in),
    .denconfig1_den_drv_cfg_rly4_out(denconfig1_den_drv_cfg_rly4_out),
    // DenConfig1.DEN_RLY_CFG_RLY4
    .denconfig1_den_rly_cfg_rly4_en(denconfig1_den_rly_cfg_rly4_en),
    .denconfig1_den_rly_cfg_rly4_in(denconfig1_den_rly_cfg_rly4_in),
    .denconfig1_den_rly_cfg_rly4_out(denconfig1_den_rly_cfg_rly4_out),

    // DenConfig2.DEN_DRV_CFG_RLY5
    .denconfig2_den_drv_cfg_rly5_en(denconfig2_den_drv_cfg_rly5_en),
    .denconfig2_den_drv_cfg_rly5_in(denconfig2_den_drv_cfg_rly5_in),
    .denconfig2_den_drv_cfg_rly5_out(denconfig2_den_drv_cfg_rly5_out),
    // DenConfig2.DEN_RLY_CFG_RLY5
    .denconfig2_den_rly_cfg_rly5_en(denconfig2_den_rly_cfg_rly5_en),
    .denconfig2_den_rly_cfg_rly5_in(denconfig2_den_rly_cfg_rly5_in),
    .denconfig2_den_rly_cfg_rly5_out(denconfig2_den_rly_cfg_rly5_out),
    // DenConfig2.DEN_DRV_CFG_RLY6
    .denconfig2_den_drv_cfg_rly6_en(denconfig2_den_drv_cfg_rly6_en),
    .denconfig2_den_drv_cfg_rly6_in(denconfig2_den_drv_cfg_rly6_in),
    .denconfig2_den_drv_cfg_rly6_out(denconfig2_den_drv_cfg_rly6_out),
    // DenConfig2.DEN_RLY_CFG_RLY6
    .denconfig2_den_rly_cfg_rly6_en(denconfig2_den_rly_cfg_rly6_en),
    .denconfig2_den_rly_cfg_rly6_in(denconfig2_den_rly_cfg_rly6_in),
    .denconfig2_den_rly_cfg_rly6_out(denconfig2_den_rly_cfg_rly6_out),
    // DenConfig2.DEN_DRV_CFG_RLY7
    .denconfig2_den_drv_cfg_rly7_en(denconfig2_den_drv_cfg_rly7_en),
    .denconfig2_den_drv_cfg_rly7_in(denconfig2_den_drv_cfg_rly7_in),
    .denconfig2_den_drv_cfg_rly7_out(denconfig2_den_drv_cfg_rly7_out),
    // DenConfig2.DEN_RLY_CFG_RLY7
    .denconfig2_den_rly_cfg_rly7_en(denconfig2_den_rly_cfg_rly7_en),
    .denconfig2_den_rly_cfg_rly7_in(denconfig2_den_rly_cfg_rly7_in),
    .denconfig2_den_rly_cfg_rly7_out(denconfig2_den_rly_cfg_rly7_out),
    // DenConfig2.DEN_DRV_CFG_RLY8
    .denconfig2_den_drv_cfg_rly8_en(denconfig2_den_drv_cfg_rly8_en),
    .denconfig2_den_drv_cfg_rly8_in(denconfig2_den_drv_cfg_rly8_in),
    .denconfig2_den_drv_cfg_rly8_out(denconfig2_den_drv_cfg_rly8_out),
    // DenConfig2.DEN_RLY_CFG_RLY8
    .denconfig2_den_rly_cfg_rly8_en(denconfig2_den_rly_cfg_rly8_en),
    .denconfig2_den_rly_cfg_rly8_in(denconfig2_den_rly_cfg_rly8_in),
    .denconfig2_den_rly_cfg_rly8_out(denconfig2_den_rly_cfg_rly8_out),

    // DenConfig3.DEN_DRV_CFG_RLY9
    .denconfig3_den_drv_cfg_rly9_en(denconfig3_den_drv_cfg_rly9_en),
    .denconfig3_den_drv_cfg_rly9_in(denconfig3_den_drv_cfg_rly9_in),
    .denconfig3_den_drv_cfg_rly9_out(denconfig3_den_drv_cfg_rly9_out),
    // DenConfig3.DEN_RLY_CFG_RLY9
    .denconfig3_den_rly_cfg_rly9_en(denconfig3_den_rly_cfg_rly9_en),
    .denconfig3_den_rly_cfg_rly9_in(denconfig3_den_rly_cfg_rly9_in),
    .denconfig3_den_rly_cfg_rly9_out(denconfig3_den_rly_cfg_rly9_out),
    // DenConfig3.DEN_DRV_CFG_VLV1
    .denconfig3_den_drv_cfg_vlv1_en(denconfig3_den_drv_cfg_vlv1_en),
    .denconfig3_den_drv_cfg_vlv1_in(denconfig3_den_drv_cfg_vlv1_in),
    .denconfig3_den_drv_cfg_vlv1_out(denconfig3_den_drv_cfg_vlv1_out),
    // DenConfig3.DEN_RLY_CFG_VLV1
    .denconfig3_den_rly_cfg_vlv1_en(denconfig3_den_rly_cfg_vlv1_en),
    .denconfig3_den_rly_cfg_vlv1_in(denconfig3_den_rly_cfg_vlv1_in),
    .denconfig3_den_rly_cfg_vlv1_out(denconfig3_den_rly_cfg_vlv1_out),
    // DenConfig3.DEN_DRV_CFG_VLV2
    .denconfig3_den_drv_cfg_vlv2_en(denconfig3_den_drv_cfg_vlv2_en),
    .denconfig3_den_drv_cfg_vlv2_in(denconfig3_den_drv_cfg_vlv2_in),
    .denconfig3_den_drv_cfg_vlv2_out(denconfig3_den_drv_cfg_vlv2_out),
    // DenConfig3.DEN_RLY_CFG_VLV2
    .denconfig3_den_rly_cfg_vlv2_en(denconfig3_den_rly_cfg_vlv2_en),
    .denconfig3_den_rly_cfg_vlv2_in(denconfig3_den_rly_cfg_vlv2_in),
    .denconfig3_den_rly_cfg_vlv2_out(denconfig3_den_rly_cfg_vlv2_out),
    // DenConfig3.DEN_DRV_CFG_VLV3
    .denconfig3_den_drv_cfg_vlv3_en(denconfig3_den_drv_cfg_vlv3_en),
    .denconfig3_den_drv_cfg_vlv3_in(denconfig3_den_drv_cfg_vlv3_in),
    .denconfig3_den_drv_cfg_vlv3_out(denconfig3_den_drv_cfg_vlv3_out),
    // DenConfig3.DEN_RLY_CFG_VLV3
    .denconfig3_den_rly_cfg_vlv3_en(denconfig3_den_rly_cfg_vlv3_en),
    .denconfig3_den_rly_cfg_vlv3_in(denconfig3_den_rly_cfg_vlv3_in),
    .denconfig3_den_rly_cfg_vlv3_out(denconfig3_den_rly_cfg_vlv3_out),

    // DenConfig4.DEN_DRV_CFG_HTR1
    .denconfig4_den_drv_cfg_htr1_en(denconfig4_den_drv_cfg_htr1_en),
    .denconfig4_den_drv_cfg_htr1_in(denconfig4_den_drv_cfg_htr1_in),
    .denconfig4_den_drv_cfg_htr1_out(denconfig4_den_drv_cfg_htr1_out),
    // DenConfig4.DEN_RLY_CFG_HTR1
    .denconfig4_den_rly_cfg_htr1_en(denconfig4_den_rly_cfg_htr1_en),
    .denconfig4_den_rly_cfg_htr1_in(denconfig4_den_rly_cfg_htr1_in),
    .denconfig4_den_rly_cfg_htr1_out(denconfig4_den_rly_cfg_htr1_out),
    // DenConfig4.DEN_DRV_CFG_HTR2
    .denconfig4_den_drv_cfg_htr2_en(denconfig4_den_drv_cfg_htr2_en),
    .denconfig4_den_drv_cfg_htr2_in(denconfig4_den_drv_cfg_htr2_in),
    .denconfig4_den_drv_cfg_htr2_out(denconfig4_den_drv_cfg_htr2_out),
    // DenConfig4.DEN_RLY_CFG_HTR2
    .denconfig4_den_rly_cfg_htr2_en(denconfig4_den_rly_cfg_htr2_en),
    .denconfig4_den_rly_cfg_htr2_in(denconfig4_den_rly_cfg_htr2_in),
    .denconfig4_den_rly_cfg_htr2_out(denconfig4_den_rly_cfg_htr2_out),
    // DenConfig4.DEN_DRV_CFG_HB1
    .denconfig4_den_drv_cfg_hb1_en(denconfig4_den_drv_cfg_hb1_en),
    .denconfig4_den_drv_cfg_hb1_in(denconfig4_den_drv_cfg_hb1_in),
    .denconfig4_den_drv_cfg_hb1_out(denconfig4_den_drv_cfg_hb1_out),
    // DenConfig4.DEN_RLY_CFG_HB1
    .denconfig4_den_rly_cfg_hb1_en(denconfig4_den_rly_cfg_hb1_en),
    .denconfig4_den_rly_cfg_hb1_in(denconfig4_den_rly_cfg_hb1_in),
    .denconfig4_den_rly_cfg_hb1_out(denconfig4_den_rly_cfg_hb1_out),
    // DenConfig4.DEN_DRV_CFG_HB2
    .denconfig4_den_drv_cfg_hb2_en(denconfig4_den_drv_cfg_hb2_en),
    .denconfig4_den_drv_cfg_hb2_in(denconfig4_den_drv_cfg_hb2_in),
    .denconfig4_den_drv_cfg_hb2_out(denconfig4_den_drv_cfg_hb2_out),
    // DenConfig4.DEN_RLY_CFG_HB2
    .denconfig4_den_rly_cfg_hb2_en(denconfig4_den_rly_cfg_hb2_en),
    .denconfig4_den_rly_cfg_hb2_in(denconfig4_den_rly_cfg_hb2_in),
    .denconfig4_den_rly_cfg_hb2_out(denconfig4_den_rly_cfg_hb2_out),

    // OEConfig0.IGN_OE
    .oeconfig0_ign_oe_en(oeconfig0_ign_oe_en),
    .oeconfig0_ign_oe_in(oeconfig0_ign_oe_in),
    .oeconfig0_ign_oe_out(oeconfig0_ign_oe_out),
    // OEConfig0.INJ_OE
    .oeconfig0_inj_oe_en(oeconfig0_inj_oe_en),
    .oeconfig0_inj_oe_in(oeconfig0_inj_oe_in),
    .oeconfig0_inj_oe_out(oeconfig0_inj_oe_out),

    // OEConfig1.RLY_OE
    .oeconfig1_rly_oe_en(oeconfig1_rly_oe_en),
    .oeconfig1_rly_oe_in(oeconfig1_rly_oe_in),
    .oeconfig1_rly_oe_out(oeconfig1_rly_oe_out),

    // OEConfig2.RLY_OE
    .oeconfig2_rly_oe_en(oeconfig2_rly_oe_en),
    .oeconfig2_rly_oe_in(oeconfig2_rly_oe_in),
    .oeconfig2_rly_oe_out(oeconfig2_rly_oe_out),
    // OEConfig2.HTR_OE
    .oeconfig2_htr_oe_en(oeconfig2_htr_oe_en),
    .oeconfig2_htr_oe_in(oeconfig2_htr_oe_in),
    .oeconfig2_htr_oe_out(oeconfig2_htr_oe_out),
    // OEConfig2.VLV_OE
    .oeconfig2_vlv_oe_en(oeconfig2_vlv_oe_en),
    .oeconfig2_vlv_oe_in(oeconfig2_vlv_oe_in),
    .oeconfig2_vlv_oe_out(oeconfig2_vlv_oe_out),

    // OEConfig3.HS_OE
    .oeconfig3_hs_oe_en(oeconfig3_hs_oe_en),
    .oeconfig3_hs_oe_in(oeconfig3_hs_oe_in),
    .oeconfig3_hs_oe_out(oeconfig3_hs_oe_out),
    // OEConfig3.LS_OE
    .oeconfig3_ls_oe_en(oeconfig3_ls_oe_en),
    .oeconfig3_ls_oe_in(oeconfig3_ls_oe_in),
    .oeconfig3_ls_oe_out(oeconfig3_ls_oe_out),

    // DDConfig0.IGN_DD
    .ddconfig0_ign_dd_en(ddconfig0_ign_dd_en),
    .ddconfig0_ign_dd_in(ddconfig0_ign_dd_in),
    .ddconfig0_ign_dd_out(ddconfig0_ign_dd_out),
    // DDConfig0.INJ_DD
    .ddconfig0_inj_dd_en(ddconfig0_inj_dd_en),
    .ddconfig0_inj_dd_in(ddconfig0_inj_dd_in),
    .ddconfig0_inj_dd_out(ddconfig0_inj_dd_out),

    // DDConfig1.RLY_DD
    .ddconfig1_rly_dd_en(ddconfig1_rly_dd_en),
    .ddconfig1_rly_dd_in(ddconfig1_rly_dd_in),
    .ddconfig1_rly_dd_out(ddconfig1_rly_dd_out),

    // DDConfig2.RLY_DD
    .ddconfig2_rly_dd_en(ddconfig2_rly_dd_en),
    .ddconfig2_rly_dd_in(ddconfig2_rly_dd_in),
    .ddconfig2_rly_dd_out(ddconfig2_rly_dd_out),
    // DDConfig2.HTR_DD
    .ddconfig2_htr_dd_en(ddconfig2_htr_dd_en),
    .ddconfig2_htr_dd_in(ddconfig2_htr_dd_in),
    .ddconfig2_htr_dd_out(ddconfig2_htr_dd_out),
    // DDConfig2.VLV_DD
    .ddconfig2_vlv_dd_en(ddconfig2_vlv_dd_en),
    .ddconfig2_vlv_dd_in(ddconfig2_vlv_dd_in),
    .ddconfig2_vlv_dd_out(ddconfig2_vlv_dd_out),
    // DDConfig2.HB_DD
    .ddconfig2_hb_dd_en(ddconfig2_hb_dd_en),
    .ddconfig2_hb_dd_in(ddconfig2_hb_dd_in),
    .ddconfig2_hb_dd_out(ddconfig2_hb_dd_out),

    // Cont0.IGN_ON
    .cont0_ign_on_en(cont0_ign_on_en),
    .cont0_ign_on_in(cont0_ign_on_in),
    .cont0_ign_on_out(cont0_ign_on_out),
    // Cont0.INJ_ON
    .cont0_inj_on_en(cont0_inj_on_en),
    .cont0_inj_on_in(cont0_inj_on_in),
    .cont0_inj_on_out(cont0_inj_on_out),

    // Cont1.RLY_ON
    .cont1_rly_on_en(cont1_rly_on_en),
    .cont1_rly_on_in(cont1_rly_on_in),
    .cont1_rly_on_out(cont1_rly_on_out),

    // Cont2.RLY_ON
    .cont2_rly_on_en(cont2_rly_on_en),
    .cont2_rly_on_in(cont2_rly_on_in),
    .cont2_rly_on_out(cont2_rly_on_out),
    // Cont2.HTR_ON
    .cont2_htr_on_en(cont2_htr_on_en),
    .cont2_htr_on_in(cont2_htr_on_in),
    .cont2_htr_on_out(cont2_htr_on_out),
    // Cont2.VLV_ON
    .cont2_vlv_on_en(cont2_vlv_on_en),
    .cont2_vlv_on_in(cont2_vlv_on_in),
    .cont2_vlv_on_out(cont2_vlv_on_out),
    // Cont2.HB_ON
    .cont2_hb_on_en(cont2_hb_on_en),
    .cont2_hb_on_in(cont2_hb_on_in),
    .cont2_hb_on_out(cont2_hb_on_out),

    // BRIConfig0.FW_MODE
    .briconfig0_fw_mode_en(briconfig0_fw_mode_en),
    .briconfig0_fw_mode_in(briconfig0_fw_mode_in),
    .briconfig0_fw_mode_out(briconfig0_fw_mode_out),
    // BRIConfig0.HS_LS_MODE
    .briconfig0_hs_ls_mode_en(briconfig0_hs_ls_mode_en),
    .briconfig0_hs_ls_mode_in(briconfig0_hs_ls_mode_in),
    .briconfig0_hs_ls_mode_out(briconfig0_hs_ls_mode_out),

    // IgnDiagConfig.EN_DIAG_OL_IGN
    .igndiagconfig_en_diag_ol_ign_en(igndiagconfig_en_diag_ol_ign_en),
    .igndiagconfig_en_diag_ol_ign_in(igndiagconfig_en_diag_ol_ign_in),
    .igndiagconfig_en_diag_ol_ign_out(igndiagconfig_en_diag_ol_ign_out),
    // IgnDiagConfig.SEL_OL_TH_IGN
    .igndiagconfig_sel_ol_th_ign_en(igndiagconfig_sel_ol_th_ign_en),
    .igndiagconfig_sel_ol_th_ign_in(igndiagconfig_sel_ol_th_ign_in),
    .igndiagconfig_sel_ol_th_ign_out(igndiagconfig_sel_ol_th_ign_out),

    // OutDiagConfig0.DIAG_INJ1
    .outdiagconfig0_diag_inj1_en(outdiagconfig0_diag_inj1_en),
    .outdiagconfig0_diag_inj1_in(outdiagconfig0_diag_inj1_in),
    .outdiagconfig0_diag_inj1_out(outdiagconfig0_diag_inj1_out),
    // OutDiagConfig0.DIAG_INJ2
    .outdiagconfig0_diag_inj2_en(outdiagconfig0_diag_inj2_en),
    .outdiagconfig0_diag_inj2_in(outdiagconfig0_diag_inj2_in),
    .outdiagconfig0_diag_inj2_out(outdiagconfig0_diag_inj2_out),
    // OutDiagConfig0.DIAG_INJ3
    .outdiagconfig0_diag_inj3_en(outdiagconfig0_diag_inj3_en),
    .outdiagconfig0_diag_inj3_in(outdiagconfig0_diag_inj3_in),
    .outdiagconfig0_diag_inj3_out(outdiagconfig0_diag_inj3_out),
    // OutDiagConfig0.DIAG_INJ4
    .outdiagconfig0_diag_inj4_en(outdiagconfig0_diag_inj4_en),
    .outdiagconfig0_diag_inj4_in(outdiagconfig0_diag_inj4_in),
    .outdiagconfig0_diag_inj4_out(outdiagconfig0_diag_inj4_out),

    // OutDiagConfig1.DIAG_RLY1
    .outdiagconfig1_diag_rly1_en(outdiagconfig1_diag_rly1_en),
    .outdiagconfig1_diag_rly1_in(outdiagconfig1_diag_rly1_in),
    .outdiagconfig1_diag_rly1_out(outdiagconfig1_diag_rly1_out),
    // OutDiagConfig1.DIAG_RLY2
    .outdiagconfig1_diag_rly2_en(outdiagconfig1_diag_rly2_en),
    .outdiagconfig1_diag_rly2_in(outdiagconfig1_diag_rly2_in),
    .outdiagconfig1_diag_rly2_out(outdiagconfig1_diag_rly2_out),
    // OutDiagConfig1.DIAG_RLY3
    .outdiagconfig1_diag_rly3_en(outdiagconfig1_diag_rly3_en),
    .outdiagconfig1_diag_rly3_in(outdiagconfig1_diag_rly3_in),
    .outdiagconfig1_diag_rly3_out(outdiagconfig1_diag_rly3_out),
    // OutDiagConfig1.DIAG_RLY4
    .outdiagconfig1_diag_rly4_en(outdiagconfig1_diag_rly4_en),
    .outdiagconfig1_diag_rly4_in(outdiagconfig1_diag_rly4_in),
    .outdiagconfig1_diag_rly4_out(outdiagconfig1_diag_rly4_out),

    // OutDiagConfig2.DIAG_RLY5
    .outdiagconfig2_diag_rly5_en(outdiagconfig2_diag_rly5_en),
    .outdiagconfig2_diag_rly5_in(outdiagconfig2_diag_rly5_in),
    .outdiagconfig2_diag_rly5_out(outdiagconfig2_diag_rly5_out),
    // OutDiagConfig2.DIAG_RLY6
    .outdiagconfig2_diag_rly6_en(outdiagconfig2_diag_rly6_en),
    .outdiagconfig2_diag_rly6_in(outdiagconfig2_diag_rly6_in),
    .outdiagconfig2_diag_rly6_out(outdiagconfig2_diag_rly6_out),
    // OutDiagConfig2.DIAG_RLY7
    .outdiagconfig2_diag_rly7_en(outdiagconfig2_diag_rly7_en),
    .outdiagconfig2_diag_rly7_in(outdiagconfig2_diag_rly7_in),
    .outdiagconfig2_diag_rly7_out(outdiagconfig2_diag_rly7_out),
    // OutDiagConfig2.DIAG_RLY8
    .outdiagconfig2_diag_rly8_en(outdiagconfig2_diag_rly8_en),
    .outdiagconfig2_diag_rly8_in(outdiagconfig2_diag_rly8_in),
    .outdiagconfig2_diag_rly8_out(outdiagconfig2_diag_rly8_out),

    // OutDiagConfig3.DIAG_RLY9
    .outdiagconfig3_diag_rly9_en(outdiagconfig3_diag_rly9_en),
    .outdiagconfig3_diag_rly9_in(outdiagconfig3_diag_rly9_in),
    .outdiagconfig3_diag_rly9_out(outdiagconfig3_diag_rly9_out),
    // OutDiagConfig3.DIAG_VLV1
    .outdiagconfig3_diag_vlv1_en(outdiagconfig3_diag_vlv1_en),
    .outdiagconfig3_diag_vlv1_in(outdiagconfig3_diag_vlv1_in),
    .outdiagconfig3_diag_vlv1_out(outdiagconfig3_diag_vlv1_out),
    // OutDiagConfig3.DIAG_VLV2
    .outdiagconfig3_diag_vlv2_en(outdiagconfig3_diag_vlv2_en),
    .outdiagconfig3_diag_vlv2_in(outdiagconfig3_diag_vlv2_in),
    .outdiagconfig3_diag_vlv2_out(outdiagconfig3_diag_vlv2_out),
    // OutDiagConfig3.DIAG_VLV3
    .outdiagconfig3_diag_vlv3_en(outdiagconfig3_diag_vlv3_en),
    .outdiagconfig3_diag_vlv3_in(outdiagconfig3_diag_vlv3_in),
    .outdiagconfig3_diag_vlv3_out(outdiagconfig3_diag_vlv3_out),

    // OutDiagConfig4.DIAG_HTR1
    .outdiagconfig4_diag_htr1_en(outdiagconfig4_diag_htr1_en),
    .outdiagconfig4_diag_htr1_in(outdiagconfig4_diag_htr1_in),
    .outdiagconfig4_diag_htr1_out(outdiagconfig4_diag_htr1_out),
    // OutDiagConfig4.DIAG_HTR2
    .outdiagconfig4_diag_htr2_en(outdiagconfig4_diag_htr2_en),
    .outdiagconfig4_diag_htr2_in(outdiagconfig4_diag_htr2_in),
    .outdiagconfig4_diag_htr2_out(outdiagconfig4_diag_htr2_out),
    // OutDiagConfig4.DIAG_HB1
    .outdiagconfig4_diag_hb1_en(outdiagconfig4_diag_hb1_en),
    .outdiagconfig4_diag_hb1_in(outdiagconfig4_diag_hb1_in),
    .outdiagconfig4_diag_hb1_out(outdiagconfig4_diag_hb1_out),
    // OutDiagConfig4.DIAG_HB2
    .outdiagconfig4_diag_hb2_en(outdiagconfig4_diag_hb2_en),
    .outdiagconfig4_diag_hb2_in(outdiagconfig4_diag_hb2_in),
    .outdiagconfig4_diag_hb2_out(outdiagconfig4_diag_hb2_out),

    // CurrLimConfig0.CURR_LIM_INJ
    .currlimconfig0_curr_lim_inj_en(currlimconfig0_curr_lim_inj_en),
    .currlimconfig0_curr_lim_inj_in(currlimconfig0_curr_lim_inj_in),
    .currlimconfig0_curr_lim_inj_out(currlimconfig0_curr_lim_inj_out),

    // CurrLimConfig1.CURR_LIM_RLY
    .currlimconfig1_curr_lim_rly_en(currlimconfig1_curr_lim_rly_en),
    .currlimconfig1_curr_lim_rly_in(currlimconfig1_curr_lim_rly_in),
    .currlimconfig1_curr_lim_rly_out(currlimconfig1_curr_lim_rly_out),

    // CurrLimConfig2.CURR_LIM_RLY
    .currlimconfig2_curr_lim_rly_en(currlimconfig2_curr_lim_rly_en),
    .currlimconfig2_curr_lim_rly_in(currlimconfig2_curr_lim_rly_in),
    .currlimconfig2_curr_lim_rly_out(currlimconfig2_curr_lim_rly_out),
    // CurrLimConfig2.CURR_LIM_VLV
    .currlimconfig2_curr_lim_vlv_en(currlimconfig2_curr_lim_vlv_en),
    .currlimconfig2_curr_lim_vlv_in(currlimconfig2_curr_lim_vlv_in),
    .currlimconfig2_curr_lim_vlv_out(currlimconfig2_curr_lim_vlv_out),
    // CurrLimConfig2.CURR_LIM_HTR
    .currlimconfig2_curr_lim_htr_en(currlimconfig2_curr_lim_htr_en),
    .currlimconfig2_curr_lim_htr_in(currlimconfig2_curr_lim_htr_in),
    .currlimconfig2_curr_lim_htr_out(currlimconfig2_curr_lim_htr_out),
    // CurrLimConfig2.CURR_LIM_HB
    .currlimconfig2_curr_lim_hb_en(currlimconfig2_curr_lim_hb_en),
    .currlimconfig2_curr_lim_hb_in(currlimconfig2_curr_lim_hb_in),
    .currlimconfig2_curr_lim_hb_out(currlimconfig2_curr_lim_hb_out),

    // DlyOffConfig.DEL_OFF_RLY
    .dlyoffconfig_del_off_rly_en(dlyoffconfig_del_off_rly_en),
    .dlyoffconfig_del_off_rly_in(dlyoffconfig_del_off_rly_in),
    .dlyoffconfig_del_off_rly_out(dlyoffconfig_del_off_rly_out),
    // DlyOffConfig.DEL_OFF_HB
    .dlyoffconfig_del_off_hb_en(dlyoffconfig_del_off_hb_en),
    .dlyoffconfig_del_off_hb_in(dlyoffconfig_del_off_hb_in),
    .dlyoffconfig_del_off_hb_out(dlyoffconfig_del_off_hb_out),

    // DinConfig0.INJ_IN1
    .dinconfig0_inj_in1_en(dinconfig0_inj_in1_en),
    .dinconfig0_inj_in1_in(dinconfig0_inj_in1_in),
    .dinconfig0_inj_in1_out(dinconfig0_inj_in1_out),
    // DinConfig0.INJ_IN2
    .dinconfig0_inj_in2_en(dinconfig0_inj_in2_en),
    .dinconfig0_inj_in2_in(dinconfig0_inj_in2_in),
    .dinconfig0_inj_in2_out(dinconfig0_inj_in2_out),

    // DinConfig1.INJ_IN3
    .dinconfig1_inj_in3_en(dinconfig1_inj_in3_en),
    .dinconfig1_inj_in3_in(dinconfig1_inj_in3_in),
    .dinconfig1_inj_in3_out(dinconfig1_inj_in3_out),
    // DinConfig1.INJ_IN4
    .dinconfig1_inj_in4_en(dinconfig1_inj_in4_en),
    .dinconfig1_inj_in4_in(dinconfig1_inj_in4_in),
    .dinconfig1_inj_in4_out(dinconfig1_inj_in4_out),

    // DinConfig2.IGN_IN1
    .dinconfig2_ign_in1_en(dinconfig2_ign_in1_en),
    .dinconfig2_ign_in1_in(dinconfig2_ign_in1_in),
    .dinconfig2_ign_in1_out(dinconfig2_ign_in1_out),
    // DinConfig2.IGN_IN2
    .dinconfig2_ign_in2_en(dinconfig2_ign_in2_en),
    .dinconfig2_ign_in2_in(dinconfig2_ign_in2_in),
    .dinconfig2_ign_in2_out(dinconfig2_ign_in2_out),

    // DinConfig3.IGN_IN3
    .dinconfig3_ign_in3_en(dinconfig3_ign_in3_en),
    .dinconfig3_ign_in3_in(dinconfig3_ign_in3_in),
    .dinconfig3_ign_in3_out(dinconfig3_ign_in3_out),
    // DinConfig3.IGN_IN4
    .dinconfig3_ign_in4_en(dinconfig3_ign_in4_en),
    .dinconfig3_ign_in4_in(dinconfig3_ign_in4_in),
    .dinconfig3_ign_in4_out(dinconfig3_ign_in4_out),

    // DinConfig4.HTR_IN1
    .dinconfig4_htr_in1_en(dinconfig4_htr_in1_en),
    .dinconfig4_htr_in1_in(dinconfig4_htr_in1_in),
    .dinconfig4_htr_in1_out(dinconfig4_htr_in1_out),
    // DinConfig4.HTR_IN2
    .dinconfig4_htr_in2_en(dinconfig4_htr_in2_en),
    .dinconfig4_htr_in2_in(dinconfig4_htr_in2_in),
    .dinconfig4_htr_in2_out(dinconfig4_htr_in2_out),

    // DinConfig5.HB_IN1
    .dinconfig5_hb_in1_en(dinconfig5_hb_in1_en),
    .dinconfig5_hb_in1_in(dinconfig5_hb_in1_in),
    .dinconfig5_hb_in1_out(dinconfig5_hb_in1_out),
    // DinConfig5.HB_IN2
    .dinconfig5_hb_in2_en(dinconfig5_hb_in2_en),
    .dinconfig5_hb_in2_in(dinconfig5_hb_in2_in),
    .dinconfig5_hb_in2_out(dinconfig5_hb_in2_out),

    // DinConfig6.RLY_IN1
    .dinconfig6_rly_in1_en(dinconfig6_rly_in1_en),
    .dinconfig6_rly_in1_in(dinconfig6_rly_in1_in),
    .dinconfig6_rly_in1_out(dinconfig6_rly_in1_out),
    // DinConfig6.RLY_IN2
    .dinconfig6_rly_in2_en(dinconfig6_rly_in2_en),
    .dinconfig6_rly_in2_in(dinconfig6_rly_in2_in),
    .dinconfig6_rly_in2_out(dinconfig6_rly_in2_out),

    // DinConfig7.RLY_IN3
    .dinconfig7_rly_in3_en(dinconfig7_rly_in3_en),
    .dinconfig7_rly_in3_in(dinconfig7_rly_in3_in),
    .dinconfig7_rly_in3_out(dinconfig7_rly_in3_out),
    // DinConfig7.RLY_IN4
    .dinconfig7_rly_in4_en(dinconfig7_rly_in4_en),
    .dinconfig7_rly_in4_in(dinconfig7_rly_in4_in),
    .dinconfig7_rly_in4_out(dinconfig7_rly_in4_out),

    // DinConfig8.RLY_IN5
    .dinconfig8_rly_in5_en(dinconfig8_rly_in5_en),
    .dinconfig8_rly_in5_in(dinconfig8_rly_in5_in),
    .dinconfig8_rly_in5_out(dinconfig8_rly_in5_out),
    // DinConfig8.RLY_IN6
    .dinconfig8_rly_in6_en(dinconfig8_rly_in6_en),
    .dinconfig8_rly_in6_in(dinconfig8_rly_in6_in),
    .dinconfig8_rly_in6_out(dinconfig8_rly_in6_out),

    // DinConfig9.RLY_IN7
    .dinconfig9_rly_in7_en(dinconfig9_rly_in7_en),
    .dinconfig9_rly_in7_in(dinconfig9_rly_in7_in),
    .dinconfig9_rly_in7_out(dinconfig9_rly_in7_out),
    // DinConfig9.RLY_IN8
    .dinconfig9_rly_in8_en(dinconfig9_rly_in8_en),
    .dinconfig9_rly_in8_in(dinconfig9_rly_in8_in),
    .dinconfig9_rly_in8_out(dinconfig9_rly_in8_out),

    // DinConfig10.RLY_IN9
    .dinconfig10_rly_in9_en(dinconfig10_rly_in9_en),
    .dinconfig10_rly_in9_in(dinconfig10_rly_in9_in),
    .dinconfig10_rly_in9_out(dinconfig10_rly_in9_out),
    // DinConfig10.VLV_IN1
    .dinconfig10_vlv_in1_en(dinconfig10_vlv_in1_en),
    .dinconfig10_vlv_in1_in(dinconfig10_vlv_in1_in),
    .dinconfig10_vlv_in1_out(dinconfig10_vlv_in1_out),

    // DinConfig11.VLV_IN2
    .dinconfig11_vlv_in2_en(dinconfig11_vlv_in2_en),
    .dinconfig11_vlv_in2_in(dinconfig11_vlv_in2_in),
    .dinconfig11_vlv_in2_out(dinconfig11_vlv_in2_out),
    // DinConfig11.VLV_IN3
    .dinconfig11_vlv_in3_en(dinconfig11_vlv_in3_en),
    .dinconfig11_vlv_in3_in(dinconfig11_vlv_in3_in),
    .dinconfig11_vlv_in3_out(dinconfig11_vlv_in3_out),

    // WDConfig0.WD_DURATION
    .wdconfig0_wd_duration_en(wdconfig0_wd_duration_en),
    .wdconfig0_wd_duration_in(wdconfig0_wd_duration_in),
    .wdconfig0_wd_duration_out(wdconfig0_wd_duration_out),
    // WDConfig0.VRS_WD_DURATION
    .wdconfig0_vrs_wd_duration_en(wdconfig0_vrs_wd_duration_en),
    .wdconfig0_vrs_wd_duration_in(wdconfig0_vrs_wd_duration_in),
    .wdconfig0_vrs_wd_duration_out(wdconfig0_vrs_wd_duration_out),
    // WDConfig0.VRS_WD_EN
    .wdconfig0_vrs_wd_en_en(wdconfig0_vrs_wd_en_en),
    .wdconfig0_vrs_wd_en_in(wdconfig0_vrs_wd_en_in),
    .wdconfig0_vrs_wd_en_out(wdconfig0_vrs_wd_en_out),

    // WDConfig1.SPI_ERR_CNT_CFG
    .wdconfig1_spi_err_cnt_cfg_en(wdconfig1_spi_err_cnt_cfg_en),
    .wdconfig1_spi_err_cnt_cfg_in(wdconfig1_spi_err_cnt_cfg_in),
    .wdconfig1_spi_err_cnt_cfg_out(wdconfig1_spi_err_cnt_cfg_out),
    // WDConfig1.SPI_RFH_CNT_CFG
    .wdconfig1_spi_rfh_cnt_cfg_en(wdconfig1_spi_rfh_cnt_cfg_en),
    .wdconfig1_spi_rfh_cnt_cfg_in(wdconfig1_spi_rfh_cnt_cfg_in),
    .wdconfig1_spi_rfh_cnt_cfg_out(wdconfig1_spi_rfh_cnt_cfg_out),
    // WDConfig1.SPI_RST_ERR_FS
    .wdconfig1_spi_rst_err_fs_en(wdconfig1_spi_rst_err_fs_en),
    .wdconfig1_spi_rst_err_fs_in(wdconfig1_spi_rst_err_fs_in),
    .wdconfig1_spi_rst_err_fs_out(wdconfig1_spi_rst_err_fs_out),

    // VrsConfig0.VRS_MODE_CFG
    .vrsconfig0_vrs_mode_cfg_en(vrsconfig0_vrs_mode_cfg_en),
    .vrsconfig0_vrs_mode_cfg_in(vrsconfig0_vrs_mode_cfg_in),
    .vrsconfig0_vrs_mode_cfg_out(vrsconfig0_vrs_mode_cfg_out),
    // VrsConfig0.VRS_REF
    .vrsconfig0_vrs_ref_en(vrsconfig0_vrs_ref_en),
    .vrsconfig0_vrs_ref_in(vrsconfig0_vrs_ref_in),
    .vrsconfig0_vrs_ref_out(vrsconfig0_vrs_ref_out),
    // VrsConfig0.VRS_TEST_CFG
    .vrsconfig0_vrs_test_cfg_en(vrsconfig0_vrs_test_cfg_en),
    .vrsconfig0_vrs_test_cfg_in(vrsconfig0_vrs_test_cfg_in),
    .vrsconfig0_vrs_test_cfg_out(vrsconfig0_vrs_test_cfg_out),
    // VrsConfig0.VRSO_SPI_CTRL_MODE
    .vrsconfig0_vrso_spi_ctrl_mode_en(vrsconfig0_vrso_spi_ctrl_mode_en),
    .vrsconfig0_vrso_spi_ctrl_mode_in(vrsconfig0_vrso_spi_ctrl_mode_in),
    .vrsconfig0_vrso_spi_ctrl_mode_out(vrsconfig0_vrso_spi_ctrl_mode_out),
    // VrsConfig0.VRSO_SPI_CTRL
    .vrsconfig0_vrso_spi_ctrl_en(vrsconfig0_vrso_spi_ctrl_en),
    .vrsconfig0_vrso_spi_ctrl_in(vrsconfig0_vrso_spi_ctrl_in),
    .vrsconfig0_vrso_spi_ctrl_out(vrsconfig0_vrso_spi_ctrl_out),

    // VrsConfig1.VRSF
    .vrsconfig1_vrsf_en(vrsconfig1_vrsf_en),
    .vrsconfig1_vrsf_in(vrsconfig1_vrsf_in),
    .vrsconfig1_vrsf_out(vrsconfig1_vrsf_out),
    // VrsConfig1.VRSM
    .vrsconfig1_vrsm_en(vrsconfig1_vrsm_en),
    .vrsconfig1_vrsm_in(vrsconfig1_vrsm_in),
    .vrsconfig1_vrsm_out(vrsconfig1_vrsm_out),
    // VrsConfig1.VRSRF
    .vrsconfig1_vrsrf_en(vrsconfig1_vrsrf_en),
    .vrsconfig1_vrsrf_in(vrsconfig1_vrsrf_in),
    .vrsconfig1_vrsrf_out(vrsconfig1_vrsrf_out),
    // VrsConfig1.VRSFF
    .vrsconfig1_vrsff_en(vrsconfig1_vrsff_en),
    .vrsconfig1_vrsff_in(vrsconfig1_vrsff_in),
    .vrsconfig1_vrsff_out(vrsconfig1_vrsff_out),
    // VrsConfig1.VRSEFF
    .vrsconfig1_vrseff_en(vrsconfig1_vrseff_en),
    .vrsconfig1_vrseff_in(vrsconfig1_vrseff_in),
    .vrsconfig1_vrseff_out(vrsconfig1_vrseff_out),
    // VrsConfig1.VRSO_EN
    .vrsconfig1_vrso_en_en(vrsconfig1_vrso_en_en),
    .vrsconfig1_vrso_en_in(vrsconfig1_vrso_en_in),
    .vrsconfig1_vrso_en_out(vrsconfig1_vrso_en_out),

    // VrsConfig2.VRS_OL_DIAG
    .vrsconfig2_vrs_ol_diag_en(vrsconfig2_vrs_ol_diag_en),
    .vrsconfig2_vrs_ol_diag_in(vrsconfig2_vrs_ol_diag_in),
    .vrsconfig2_vrs_ol_diag_out(vrsconfig2_vrs_ol_diag_out),

    // MscConfig0.MSC_CLK_DIV_CFG
    .mscconfig0_msc_clk_div_cfg_en(mscconfig0_msc_clk_div_cfg_en),
    .mscconfig0_msc_clk_div_cfg_in(mscconfig0_msc_clk_div_cfg_in),
    .mscconfig0_msc_clk_div_cfg_out(mscconfig0_msc_clk_div_cfg_out),
    // MscConfig0.MSC_SV_EN
    .mscconfig0_msc_sv_en_en(mscconfig0_msc_sv_en_en),
    .mscconfig0_msc_sv_en_in(mscconfig0_msc_sv_en_in),
    .mscconfig0_msc_sv_en_out(mscconfig0_msc_sv_en_out),

    // MscConfig1.MSC_CRC_CFG
    .mscconfig1_msc_crc_cfg_en(mscconfig1_msc_crc_cfg_en),
    .mscconfig1_msc_crc_cfg_in(mscconfig1_msc_crc_cfg_in),
    .mscconfig1_msc_crc_cfg_out(mscconfig1_msc_crc_cfg_out),
    // MscConfig1.MSC_UP_FRAME
    .mscconfig1_msc_up_frame_en(mscconfig1_msc_up_frame_en),
    .mscconfig1_msc_up_frame_in(mscconfig1_msc_up_frame_in),
    .mscconfig1_msc_up_frame_out(mscconfig1_msc_up_frame_out),
    // MscConfig1.MSC_ADDR_MODE
    .mscconfig1_msc_addr_mode_en(mscconfig1_msc_addr_mode_en),
    .mscconfig1_msc_addr_mode_in(mscconfig1_msc_addr_mode_in),
    .mscconfig1_msc_addr_mode_out(mscconfig1_msc_addr_mode_out),
    // MscConfig1.MSC_ADDR_CFG
    .mscconfig1_msc_addr_cfg_en(mscconfig1_msc_addr_cfg_en),
    .mscconfig1_msc_addr_cfg_in(mscconfig1_msc_addr_cfg_in),
    .mscconfig1_msc_addr_cfg_out(mscconfig1_msc_addr_cfg_out),
    // MscConfig1.OD_MISO
    .mscconfig1_od_miso_en(mscconfig1_od_miso_en),
    .mscconfig1_od_miso_in(mscconfig1_od_miso_in),
    .mscconfig1_od_miso_out(mscconfig1_od_miso_out),

    // AoutConfig.AMUX
    .aoutconfig_amux_en(aoutconfig_amux_en),
    .aoutconfig_amux_in(aoutconfig_amux_in),
    .aoutconfig_amux_out(aoutconfig_amux_out),
    // AoutConfig.VDDIO_RNG
    .aoutconfig_vddio_rng_en(aoutconfig_vddio_rng_en),
    .aoutconfig_vddio_rng_in(aoutconfig_vddio_rng_in),
    .aoutconfig_vddio_rng_out(aoutconfig_vddio_rng_out),
    // AoutConfig.VPWR_RNG
    .aoutconfig_vpwr_rng_en(aoutconfig_vpwr_rng_en),
    .aoutconfig_vpwr_rng_in(aoutconfig_vpwr_rng_in),
    .aoutconfig_vpwr_rng_out(aoutconfig_vpwr_rng_out),

    // RstbConfig.VDD5_UV_RSTB_CFG
    .rstbconfig_vdd5_uv_rstb_cfg_en(rstbconfig_vdd5_uv_rstb_cfg_en),
    .rstbconfig_vdd5_uv_rstb_cfg_in(rstbconfig_vdd5_uv_rstb_cfg_in),
    .rstbconfig_vdd5_uv_rstb_cfg_out(rstbconfig_vdd5_uv_rstb_cfg_out),
    // RstbConfig.VDD5_OV_RSTB_CFG
    .rstbconfig_vdd5_ov_rstb_cfg_en(rstbconfig_vdd5_ov_rstb_cfg_en),
    .rstbconfig_vdd5_ov_rstb_cfg_in(rstbconfig_vdd5_ov_rstb_cfg_in),
    .rstbconfig_vdd5_ov_rstb_cfg_out(rstbconfig_vdd5_ov_rstb_cfg_out),
    // RstbConfig.WD_RSTB_CFG
    .rstbconfig_wd_rstb_cfg_en(rstbconfig_wd_rstb_cfg_en),
    .rstbconfig_wd_rstb_cfg_in(rstbconfig_wd_rstb_cfg_in),
    .rstbconfig_wd_rstb_cfg_out(rstbconfig_wd_rstb_cfg_out),

    // FaultbConfig0.WD_SV_FAIL_DIAG
    .faultbconfig0_wd_sv_fail_diag_en(faultbconfig0_wd_sv_fail_diag_en),
    .faultbconfig0_wd_sv_fail_diag_in(faultbconfig0_wd_sv_fail_diag_in),
    .faultbconfig0_wd_sv_fail_diag_out(faultbconfig0_wd_sv_fail_diag_out),
    // FaultbConfig0.SPI_MSC_FAIL_DIAG
    .faultbconfig0_spi_msc_fail_diag_en(faultbconfig0_spi_msc_fail_diag_en),
    .faultbconfig0_spi_msc_fail_diag_in(faultbconfig0_spi_msc_fail_diag_in),
    .faultbconfig0_spi_msc_fail_diag_out(faultbconfig0_spi_msc_fail_diag_out),
    // FaultbConfig0.OTP_FAIL_DIAG
    .faultbconfig0_otp_fail_diag_en(faultbconfig0_otp_fail_diag_en),
    .faultbconfig0_otp_fail_diag_in(faultbconfig0_otp_fail_diag_in),
    .faultbconfig0_otp_fail_diag_out(faultbconfig0_otp_fail_diag_out),
    // FaultbConfig0.FAULT_VRS_WD_DIAG
    .faultbconfig0_fault_vrs_wd_diag_en(faultbconfig0_fault_vrs_wd_diag_en),
    .faultbconfig0_fault_vrs_wd_diag_in(faultbconfig0_fault_vrs_wd_diag_in),
    .faultbconfig0_fault_vrs_wd_diag_out(faultbconfig0_fault_vrs_wd_diag_out),
    // FaultbConfig0.VRS_OL_SC_DIAG
    .faultbconfig0_vrs_ol_sc_diag_en(faultbconfig0_vrs_ol_sc_diag_en),
    .faultbconfig0_vrs_ol_sc_diag_in(faultbconfig0_vrs_ol_sc_diag_in),
    .faultbconfig0_vrs_ol_sc_diag_out(faultbconfig0_vrs_ol_sc_diag_out),
    // FaultbConfig0.GND_FAIL_DIAG
    .faultbconfig0_gnd_fail_diag_en(faultbconfig0_gnd_fail_diag_en),
    .faultbconfig0_gnd_fail_diag_in(faultbconfig0_gnd_fail_diag_in),
    .faultbconfig0_gnd_fail_diag_out(faultbconfig0_gnd_fail_diag_out),
    // FaultbConfig0.FAULTB_LATCH_DATA
    .faultbconfig0_faultb_latch_data_en(faultbconfig0_faultb_latch_data_en),
    .faultbconfig0_faultb_latch_data_in(faultbconfig0_faultb_latch_data_in),
    .faultbconfig0_faultb_latch_data_out(faultbconfig0_faultb_latch_data_out),

    // FaultbConfig1.SUP_REGL_DIAG
    .faultbconfig1_sup_regl_diag_en(faultbconfig1_sup_regl_diag_en),
    .faultbconfig1_sup_regl_diag_in(faultbconfig1_sup_regl_diag_in),
    .faultbconfig1_sup_regl_diag_out(faultbconfig1_sup_regl_diag_out),
    // FaultbConfig1.CP_UV_DIAG
    .faultbconfig1_cp_uv_diag_en(faultbconfig1_cp_uv_diag_en),
    .faultbconfig1_cp_uv_diag_in(faultbconfig1_cp_uv_diag_in),
    .faultbconfig1_cp_uv_diag_out(faultbconfig1_cp_uv_diag_out),
    // FaultbConfig1.VDDIO_UV_DIAG
    .faultbconfig1_vddio_uv_diag_en(faultbconfig1_vddio_uv_diag_en),
    .faultbconfig1_vddio_uv_diag_in(faultbconfig1_vddio_uv_diag_in),
    .faultbconfig1_vddio_uv_diag_out(faultbconfig1_vddio_uv_diag_out),
    // FaultbConfig1.VDDIO_OV_DIAG
    .faultbconfig1_vddio_ov_diag_en(faultbconfig1_vddio_ov_diag_en),
    .faultbconfig1_vddio_ov_diag_in(faultbconfig1_vddio_ov_diag_in),
    .faultbconfig1_vddio_ov_diag_out(faultbconfig1_vddio_ov_diag_out),
    // FaultbConfig1.VPWR_UV_DIAG
    .faultbconfig1_vpwr_uv_diag_en(faultbconfig1_vpwr_uv_diag_en),
    .faultbconfig1_vpwr_uv_diag_in(faultbconfig1_vpwr_uv_diag_in),
    .faultbconfig1_vpwr_uv_diag_out(faultbconfig1_vpwr_uv_diag_out),
    // FaultbConfig1.VPWR_OV_DIAG
    .faultbconfig1_vpwr_ov_diag_en(faultbconfig1_vpwr_ov_diag_en),
    .faultbconfig1_vpwr_ov_diag_in(faultbconfig1_vpwr_ov_diag_in),
    .faultbconfig1_vpwr_ov_diag_out(faultbconfig1_vpwr_ov_diag_out),
    // FaultbConfig1.VDD5_UV_DIAG
    .faultbconfig1_vdd5_uv_diag_en(faultbconfig1_vdd5_uv_diag_en),
    .faultbconfig1_vdd5_uv_diag_in(faultbconfig1_vdd5_uv_diag_in),
    .faultbconfig1_vdd5_uv_diag_out(faultbconfig1_vdd5_uv_diag_out),
    // FaultbConfig1.VDD5_OV_DIAG
    .faultbconfig1_vdd5_ov_diag_en(faultbconfig1_vdd5_ov_diag_en),
    .faultbconfig1_vdd5_ov_diag_in(faultbconfig1_vdd5_ov_diag_in),
    .faultbconfig1_vdd5_ov_diag_out(faultbconfig1_vdd5_ov_diag_out),

    // FaultbConfig2.OL_SC_DIAG
    .faultbconfig2_ol_sc_diag_en(faultbconfig2_ol_sc_diag_en),
    .faultbconfig2_ol_sc_diag_in(faultbconfig2_ol_sc_diag_in),
    .faultbconfig2_ol_sc_diag_out(faultbconfig2_ol_sc_diag_out),
    // FaultbConfig2.TSD_DIAG
    .faultbconfig2_tsd_diag_en(faultbconfig2_tsd_diag_en),
    .faultbconfig2_tsd_diag_in(faultbconfig2_tsd_diag_in),
    .faultbconfig2_tsd_diag_out(faultbconfig2_tsd_diag_out),
    // FaultbConfig2.OC_DIAG
    .faultbconfig2_oc_diag_en(faultbconfig2_oc_diag_en),
    .faultbconfig2_oc_diag_in(faultbconfig2_oc_diag_in),
    .faultbconfig2_oc_diag_out(faultbconfig2_oc_diag_out),
    // FaultbConfig2.SC_IGN_DIAG
    .faultbconfig2_sc_ign_diag_en(faultbconfig2_sc_ign_diag_en),
    .faultbconfig2_sc_ign_diag_in(faultbconfig2_sc_ign_diag_in),
    .faultbconfig2_sc_ign_diag_out(faultbconfig2_sc_ign_diag_out),
    // FaultbConfig2.OL_IGN_DIAG
    .faultbconfig2_ol_ign_diag_en(faultbconfig2_ol_ign_diag_en),
    .faultbconfig2_ol_ign_diag_in(faultbconfig2_ol_ign_diag_in),
    .faultbconfig2_ol_ign_diag_out(faultbconfig2_ol_ign_diag_out),
    // FaultbConfig2.DNDIS_DRV_DIAG
    .faultbconfig2_dndis_drv_diag_en(faultbconfig2_dndis_drv_diag_en),
    .faultbconfig2_dndis_drv_diag_in(faultbconfig2_dndis_drv_diag_in),
    .faultbconfig2_dndis_drv_diag_out(faultbconfig2_dndis_drv_diag_out),
    // FaultbConfig2.FAULTB_SPI_CTRL_MODE
    .faultbconfig2_faultb_spi_ctrl_mode_en(faultbconfig2_faultb_spi_ctrl_mode_en),
    .faultbconfig2_faultb_spi_ctrl_mode_in(faultbconfig2_faultb_spi_ctrl_mode_in),
    .faultbconfig2_faultb_spi_ctrl_mode_out(faultbconfig2_faultb_spi_ctrl_mode_out),
    // FaultbConfig2.FAULTB_SPI_CTRL
    .faultbconfig2_faultb_spi_ctrl_en(faultbconfig2_faultb_spi_ctrl_en),
    .faultbconfig2_faultb_spi_ctrl_in(faultbconfig2_faultb_spi_ctrl_in),
    .faultbconfig2_faultb_spi_ctrl_out(faultbconfig2_faultb_spi_ctrl_out),

    // VrsDiag.FAULT_VRS_WD
    .vrsdiag_fault_vrs_wd_en(vrsdiag_fault_vrs_wd_en),
    .vrsdiag_fault_vrs_wd_in(vrsdiag_fault_vrs_wd_in),
    // VrsDiag.VRS_SCB
    .vrsdiag_vrs_scb_en(vrsdiag_vrs_scb_en),
    .vrsdiag_vrs_scb_in(vrsdiag_vrs_scb_in),
    // VrsDiag.VRS_SCG
    .vrsdiag_vrs_scg_en(vrsdiag_vrs_scg_en),
    .vrsdiag_vrs_scg_in(vrsdiag_vrs_scg_in),
    // VrsDiag.VRS_OL
    .vrsdiag_vrs_ol_en(vrsdiag_vrs_ol_en),
    .vrsdiag_vrs_ol_in(vrsdiag_vrs_ol_in),
    // VrsDiag.VRS_TH_FAULT
    .vrsdiag_vrs_th_fault_en(vrsdiag_vrs_th_fault_en),
    .vrsdiag_vrs_th_fault_in(vrsdiag_vrs_th_fault_in),

    // SupDiag.SUP_REGL
    .supdiag_sup_regl_en(supdiag_sup_regl_en),
    .supdiag_sup_regl_in(supdiag_sup_regl_in),
    // SupDiag.CP_UV
    .supdiag_cp_uv_en(supdiag_cp_uv_en),
    .supdiag_cp_uv_in(supdiag_cp_uv_in),
    // SupDiag.VDDIO_UV
    .supdiag_vddio_uv_en(supdiag_vddio_uv_en),
    .supdiag_vddio_uv_in(supdiag_vddio_uv_in),
    // SupDiag.VDDIO_OV
    .supdiag_vddio_ov_en(supdiag_vddio_ov_en),
    .supdiag_vddio_ov_in(supdiag_vddio_ov_in),
    // SupDiag.VPWR_UV
    .supdiag_vpwr_uv_en(supdiag_vpwr_uv_en),
    .supdiag_vpwr_uv_in(supdiag_vpwr_uv_in),
    // SupDiag.VPWR_OV
    .supdiag_vpwr_ov_en(supdiag_vpwr_ov_en),
    .supdiag_vpwr_ov_in(supdiag_vpwr_ov_in),
    // SupDiag.VDD5_UV
    .supdiag_vdd5_uv_en(supdiag_vdd5_uv_en),
    .supdiag_vdd5_uv_in(supdiag_vdd5_uv_in),
    // SupDiag.VDD5_OV
    .supdiag_vdd5_ov_en(supdiag_vdd5_ov_en),
    .supdiag_vdd5_ov_in(supdiag_vdd5_ov_in),

    // ExtDiag0.MSC_SPI_ERROR
    .extdiag0_msc_spi_error_en(extdiag0_msc_spi_error_en),
    .extdiag0_msc_spi_error_in(extdiag0_msc_spi_error_in),
    // ExtDiag0.MSC_SV_ERROR
    .extdiag0_msc_sv_error_en(extdiag0_msc_sv_error_en),
    .extdiag0_msc_sv_error_in(extdiag0_msc_sv_error_in),
    // ExtDiag0.WD_WARN
    .extdiag0_wd_warn_en(extdiag0_wd_warn_en),
    .extdiag0_wd_warn_in(extdiag0_wd_warn_in),
    // ExtDiag0.WD_FAIL
    .extdiag0_wd_fail_en(extdiag0_wd_fail_en),
    .extdiag0_wd_fail_in(extdiag0_wd_fail_in),
    // ExtDiag0.FUSE_CHECK_ERROR
    .extdiag0_fuse_check_error_en(extdiag0_fuse_check_error_en),
    .extdiag0_fuse_check_error_in(extdiag0_fuse_check_error_in),
    // ExtDiag0.OTP_USAGE_FAULT
    .extdiag0_otp_usage_fault_en(extdiag0_otp_usage_fault_en),
    .extdiag0_otp_usage_fault_in(extdiag0_otp_usage_fault_in),
    // ExtDiag0.SELF_TEST_ERROR
    .extdiag0_self_test_error_en(extdiag0_self_test_error_en),
    .extdiag0_self_test_error_in(extdiag0_self_test_error_in),

    // ExtDiag1.PGND_LOSS
    .extdiag1_pgnd_loss_en(extdiag1_pgnd_loss_en),
    .extdiag1_pgnd_loss_in(extdiag1_pgnd_loss_in),
    // ExtDiag1.AGND_LOSS
    .extdiag1_agnd_loss_en(extdiag1_agnd_loss_en),
    .extdiag1_agnd_loss_in(extdiag1_agnd_loss_in),
    // ExtDiag1.GNDIO_LOSS
    .extdiag1_gndio_loss_en(extdiag1_gndio_loss_en),
    .extdiag1_gndio_loss_in(extdiag1_gndio_loss_in),
    // ExtDiag1.VDIG_1P5V_OV
    .extdiag1_vdig_1p5v_ov_en(extdiag1_vdig_1p5v_ov_en),
    .extdiag1_vdig_1p5v_ov_in(extdiag1_vdig_1p5v_ov_in),
    // ExtDiag1.VDIG_1P5V_UV
    .extdiag1_vdig_1p5v_uv_en(extdiag1_vdig_1p5v_uv_en),
    .extdiag1_vdig_1p5v_uv_in(extdiag1_vdig_1p5v_uv_in),
    // ExtDiag1.VANA_1P5V_UV
    .extdiag1_vana_1p5v_uv_en(extdiag1_vana_1p5v_uv_en),
    .extdiag1_vana_1p5v_uv_in(extdiag1_vana_1p5v_uv_in),
    // ExtDiag1.VANA_1P5V_OV
    .extdiag1_vana_1p5v_ov_en(extdiag1_vana_1p5v_ov_en),
    .extdiag1_vana_1p5v_ov_in(extdiag1_vana_1p5v_ov_in),
    // ExtDiag1.DIS_DRV
    .extdiag1_dis_drv_en(extdiag1_dis_drv_en),
    .extdiag1_dis_drv_in(extdiag1_dis_drv_in),

    // InjDiag0.SCG_INJ1
    .injdiag0_scg_inj1_en(injdiag0_scg_inj1_en),
    .injdiag0_scg_inj1_in(injdiag0_scg_inj1_in),
    // InjDiag0.OL_INJ1
    .injdiag0_ol_inj1_en(injdiag0_ol_inj1_en),
    .injdiag0_ol_inj1_in(injdiag0_ol_inj1_in),
    // InjDiag0.TSD_INJ1
    .injdiag0_tsd_inj1_en(injdiag0_tsd_inj1_en),
    .injdiag0_tsd_inj1_in(injdiag0_tsd_inj1_in),
    // InjDiag0.OC_INJ1
    .injdiag0_oc_inj1_en(injdiag0_oc_inj1_en),
    .injdiag0_oc_inj1_in(injdiag0_oc_inj1_in),
    // InjDiag0.SCG_INJ2
    .injdiag0_scg_inj2_en(injdiag0_scg_inj2_en),
    .injdiag0_scg_inj2_in(injdiag0_scg_inj2_in),
    // InjDiag0.OL_INJ2
    .injdiag0_ol_inj2_en(injdiag0_ol_inj2_en),
    .injdiag0_ol_inj2_in(injdiag0_ol_inj2_in),
    // InjDiag0.TSD_INJ2
    .injdiag0_tsd_inj2_en(injdiag0_tsd_inj2_en),
    .injdiag0_tsd_inj2_in(injdiag0_tsd_inj2_in),
    // InjDiag0.OC_INJ2
    .injdiag0_oc_inj2_en(injdiag0_oc_inj2_en),
    .injdiag0_oc_inj2_in(injdiag0_oc_inj2_in),

    // InjDiag1.SCG_INJ3
    .injdiag1_scg_inj3_en(injdiag1_scg_inj3_en),
    .injdiag1_scg_inj3_in(injdiag1_scg_inj3_in),
    // InjDiag1.OL_INJ3
    .injdiag1_ol_inj3_en(injdiag1_ol_inj3_en),
    .injdiag1_ol_inj3_in(injdiag1_ol_inj3_in),
    // InjDiag1.TSD_INJ3
    .injdiag1_tsd_inj3_en(injdiag1_tsd_inj3_en),
    .injdiag1_tsd_inj3_in(injdiag1_tsd_inj3_in),
    // InjDiag1.OC_INJ3
    .injdiag1_oc_inj3_en(injdiag1_oc_inj3_en),
    .injdiag1_oc_inj3_in(injdiag1_oc_inj3_in),
    // InjDiag1.SCG_INJ4
    .injdiag1_scg_inj4_en(injdiag1_scg_inj4_en),
    .injdiag1_scg_inj4_in(injdiag1_scg_inj4_in),
    // InjDiag1.OL_INJ4
    .injdiag1_ol_inj4_en(injdiag1_ol_inj4_en),
    .injdiag1_ol_inj4_in(injdiag1_ol_inj4_in),
    // InjDiag1.TSD_INJ4
    .injdiag1_tsd_inj4_en(injdiag1_tsd_inj4_en),
    .injdiag1_tsd_inj4_in(injdiag1_tsd_inj4_in),
    // InjDiag1.OC_INJ4
    .injdiag1_oc_inj4_en(injdiag1_oc_inj4_en),
    .injdiag1_oc_inj4_in(injdiag1_oc_inj4_in),

    // IgnDiag0.SCG_IGN1
    .igndiag0_scg_ign1_en(igndiag0_scg_ign1_en),
    .igndiag0_scg_ign1_in(igndiag0_scg_ign1_in),
    // IgnDiag0.OL_IGN1
    .igndiag0_ol_ign1_en(igndiag0_ol_ign1_en),
    .igndiag0_ol_ign1_in(igndiag0_ol_ign1_in),
    // IgnDiag0.SCB_IGN1
    .igndiag0_scb_ign1_en(igndiag0_scb_ign1_en),
    .igndiag0_scb_ign1_in(igndiag0_scb_ign1_in),
    // IgnDiag0.SCG_IGN2
    .igndiag0_scg_ign2_en(igndiag0_scg_ign2_en),
    .igndiag0_scg_ign2_in(igndiag0_scg_ign2_in),
    // IgnDiag0.OL_IGN2
    .igndiag0_ol_ign2_en(igndiag0_ol_ign2_en),
    .igndiag0_ol_ign2_in(igndiag0_ol_ign2_in),
    // IgnDiag0.SCB_IGN2
    .igndiag0_scb_ign2_en(igndiag0_scb_ign2_en),
    .igndiag0_scb_ign2_in(igndiag0_scb_ign2_in),
    // IgnDiag0.TSD_IGN1
    .igndiag0_tsd_ign1_en(igndiag0_tsd_ign1_en),
    .igndiag0_tsd_ign1_in(igndiag0_tsd_ign1_in),

    // IgnDiag1.SCG_IGN3
    .igndiag1_scg_ign3_en(igndiag1_scg_ign3_en),
    .igndiag1_scg_ign3_in(igndiag1_scg_ign3_in),
    // IgnDiag1.OL_IGN3
    .igndiag1_ol_ign3_en(igndiag1_ol_ign3_en),
    .igndiag1_ol_ign3_in(igndiag1_ol_ign3_in),
    // IgnDiag1.SCB_IGN3
    .igndiag1_scb_ign3_en(igndiag1_scb_ign3_en),
    .igndiag1_scb_ign3_in(igndiag1_scb_ign3_in),
    // IgnDiag1.SCG_IGN4
    .igndiag1_scg_ign4_en(igndiag1_scg_ign4_en),
    .igndiag1_scg_ign4_in(igndiag1_scg_ign4_in),
    // IgnDiag1.OL_IGN4
    .igndiag1_ol_ign4_en(igndiag1_ol_ign4_en),
    .igndiag1_ol_ign4_in(igndiag1_ol_ign4_in),
    // IgnDiag1.SCB_IGN4
    .igndiag1_scb_ign4_en(igndiag1_scb_ign4_en),
    .igndiag1_scb_ign4_in(igndiag1_scb_ign4_in),
    // IgnDiag1.TSD_IGN2
    .igndiag1_tsd_ign2_en(igndiag1_tsd_ign2_en),
    .igndiag1_tsd_ign2_in(igndiag1_tsd_ign2_in),

    // HtrDiag0.SCG_HTR1
    .htrdiag0_scg_htr1_en(htrdiag0_scg_htr1_en),
    .htrdiag0_scg_htr1_in(htrdiag0_scg_htr1_in),
    // HtrDiag0.OL_HTR1
    .htrdiag0_ol_htr1_en(htrdiag0_ol_htr1_en),
    .htrdiag0_ol_htr1_in(htrdiag0_ol_htr1_in),
    // HtrDiag0.TSD_HTR1
    .htrdiag0_tsd_htr1_en(htrdiag0_tsd_htr1_en),
    .htrdiag0_tsd_htr1_in(htrdiag0_tsd_htr1_in),
    // HtrDiag0.OC_HTR1
    .htrdiag0_oc_htr1_en(htrdiag0_oc_htr1_en),
    .htrdiag0_oc_htr1_in(htrdiag0_oc_htr1_in),
    // HtrDiag0.SCG_HTR2
    .htrdiag0_scg_htr2_en(htrdiag0_scg_htr2_en),
    .htrdiag0_scg_htr2_in(htrdiag0_scg_htr2_in),
    // HtrDiag0.OL_HTR2
    .htrdiag0_ol_htr2_en(htrdiag0_ol_htr2_en),
    .htrdiag0_ol_htr2_in(htrdiag0_ol_htr2_in),
    // HtrDiag0.TSD_HTR2
    .htrdiag0_tsd_htr2_en(htrdiag0_tsd_htr2_en),
    .htrdiag0_tsd_htr2_in(htrdiag0_tsd_htr2_in),
    // HtrDiag0.OC_HTR2
    .htrdiag0_oc_htr2_en(htrdiag0_oc_htr2_en),
    .htrdiag0_oc_htr2_in(htrdiag0_oc_htr2_in),

    // RlyDiag0.SCG_RLY1
    .rlydiag0_scg_rly1_en(rlydiag0_scg_rly1_en),
    .rlydiag0_scg_rly1_in(rlydiag0_scg_rly1_in),
    // RlyDiag0.OL_RLY1
    .rlydiag0_ol_rly1_en(rlydiag0_ol_rly1_en),
    .rlydiag0_ol_rly1_in(rlydiag0_ol_rly1_in),
    // RlyDiag0.TSD_RLY1
    .rlydiag0_tsd_rly1_en(rlydiag0_tsd_rly1_en),
    .rlydiag0_tsd_rly1_in(rlydiag0_tsd_rly1_in),
    // RlyDiag0.OC_RLY1
    .rlydiag0_oc_rly1_en(rlydiag0_oc_rly1_en),
    .rlydiag0_oc_rly1_in(rlydiag0_oc_rly1_in),
    // RlyDiag0.SCG_RLY2
    .rlydiag0_scg_rly2_en(rlydiag0_scg_rly2_en),
    .rlydiag0_scg_rly2_in(rlydiag0_scg_rly2_in),
    // RlyDiag0.OL_RLY2
    .rlydiag0_ol_rly2_en(rlydiag0_ol_rly2_en),
    .rlydiag0_ol_rly2_in(rlydiag0_ol_rly2_in),
    // RlyDiag0.TSD_RLY2
    .rlydiag0_tsd_rly2_en(rlydiag0_tsd_rly2_en),
    .rlydiag0_tsd_rly2_in(rlydiag0_tsd_rly2_in),
    // RlyDiag0.OC_RLY2
    .rlydiag0_oc_rly2_en(rlydiag0_oc_rly2_en),
    .rlydiag0_oc_rly2_in(rlydiag0_oc_rly2_in),

    // RlyDiag1.SCG_RLY3
    .rlydiag1_scg_rly3_en(rlydiag1_scg_rly3_en),
    .rlydiag1_scg_rly3_in(rlydiag1_scg_rly3_in),
    // RlyDiag1.OL_RLY3
    .rlydiag1_ol_rly3_en(rlydiag1_ol_rly3_en),
    .rlydiag1_ol_rly3_in(rlydiag1_ol_rly3_in),
    // RlyDiag1.TSD_RLY3
    .rlydiag1_tsd_rly3_en(rlydiag1_tsd_rly3_en),
    .rlydiag1_tsd_rly3_in(rlydiag1_tsd_rly3_in),
    // RlyDiag1.OC_RLY3
    .rlydiag1_oc_rly3_en(rlydiag1_oc_rly3_en),
    .rlydiag1_oc_rly3_in(rlydiag1_oc_rly3_in),
    // RlyDiag1.SCG_RLY4
    .rlydiag1_scg_rly4_en(rlydiag1_scg_rly4_en),
    .rlydiag1_scg_rly4_in(rlydiag1_scg_rly4_in),
    // RlyDiag1.OL_RLY4
    .rlydiag1_ol_rly4_en(rlydiag1_ol_rly4_en),
    .rlydiag1_ol_rly4_in(rlydiag1_ol_rly4_in),
    // RlyDiag1.TSD_RLY4
    .rlydiag1_tsd_rly4_en(rlydiag1_tsd_rly4_en),
    .rlydiag1_tsd_rly4_in(rlydiag1_tsd_rly4_in),
    // RlyDiag1.OC_RLY4
    .rlydiag1_oc_rly4_en(rlydiag1_oc_rly4_en),
    .rlydiag1_oc_rly4_in(rlydiag1_oc_rly4_in),

    // RlyDiag2.SCG_RLY5
    .rlydiag2_scg_rly5_en(rlydiag2_scg_rly5_en),
    .rlydiag2_scg_rly5_in(rlydiag2_scg_rly5_in),
    // RlyDiag2.OL_RLY5
    .rlydiag2_ol_rly5_en(rlydiag2_ol_rly5_en),
    .rlydiag2_ol_rly5_in(rlydiag2_ol_rly5_in),
    // RlyDiag2.TSD_RLY5
    .rlydiag2_tsd_rly5_en(rlydiag2_tsd_rly5_en),
    .rlydiag2_tsd_rly5_in(rlydiag2_tsd_rly5_in),
    // RlyDiag2.OC_RLY5
    .rlydiag2_oc_rly5_en(rlydiag2_oc_rly5_en),
    .rlydiag2_oc_rly5_in(rlydiag2_oc_rly5_in),
    // RlyDiag2.SCG_RLY6
    .rlydiag2_scg_rly6_en(rlydiag2_scg_rly6_en),
    .rlydiag2_scg_rly6_in(rlydiag2_scg_rly6_in),
    // RlyDiag2.OL_RLY6
    .rlydiag2_ol_rly6_en(rlydiag2_ol_rly6_en),
    .rlydiag2_ol_rly6_in(rlydiag2_ol_rly6_in),
    // RlyDiag2.TSD_RLY6
    .rlydiag2_tsd_rly6_en(rlydiag2_tsd_rly6_en),
    .rlydiag2_tsd_rly6_in(rlydiag2_tsd_rly6_in),
    // RlyDiag2.OC_RLY6
    .rlydiag2_oc_rly6_en(rlydiag2_oc_rly6_en),
    .rlydiag2_oc_rly6_in(rlydiag2_oc_rly6_in),

    // RlyDiag3.SCG_RLY7
    .rlydiag3_scg_rly7_en(rlydiag3_scg_rly7_en),
    .rlydiag3_scg_rly7_in(rlydiag3_scg_rly7_in),
    // RlyDiag3.OL_RLY7
    .rlydiag3_ol_rly7_en(rlydiag3_ol_rly7_en),
    .rlydiag3_ol_rly7_in(rlydiag3_ol_rly7_in),
    // RlyDiag3.TSD_RLY7
    .rlydiag3_tsd_rly7_en(rlydiag3_tsd_rly7_en),
    .rlydiag3_tsd_rly7_in(rlydiag3_tsd_rly7_in),
    // RlyDiag3.OC_RLY7
    .rlydiag3_oc_rly7_en(rlydiag3_oc_rly7_en),
    .rlydiag3_oc_rly7_in(rlydiag3_oc_rly7_in),
    // RlyDiag3.SCG_RLY8
    .rlydiag3_scg_rly8_en(rlydiag3_scg_rly8_en),
    .rlydiag3_scg_rly8_in(rlydiag3_scg_rly8_in),
    // RlyDiag3.OL_RLY8
    .rlydiag3_ol_rly8_en(rlydiag3_ol_rly8_en),
    .rlydiag3_ol_rly8_in(rlydiag3_ol_rly8_in),
    // RlyDiag3.TSD_RLY8
    .rlydiag3_tsd_rly8_en(rlydiag3_tsd_rly8_en),
    .rlydiag3_tsd_rly8_in(rlydiag3_tsd_rly8_in),
    // RlyDiag3.OC_RLY8
    .rlydiag3_oc_rly8_en(rlydiag3_oc_rly8_en),
    .rlydiag3_oc_rly8_in(rlydiag3_oc_rly8_in),

    // RlyDiag4.SCG_RLY9
    .rlydiag4_scg_rly9_en(rlydiag4_scg_rly9_en),
    .rlydiag4_scg_rly9_in(rlydiag4_scg_rly9_in),
    // RlyDiag4.OL_RLY9
    .rlydiag4_ol_rly9_en(rlydiag4_ol_rly9_en),
    .rlydiag4_ol_rly9_in(rlydiag4_ol_rly9_in),
    // RlyDiag4.TSD_RLY9
    .rlydiag4_tsd_rly9_en(rlydiag4_tsd_rly9_en),
    .rlydiag4_tsd_rly9_in(rlydiag4_tsd_rly9_in),
    // RlyDiag4.OC_RLY9
    .rlydiag4_oc_rly9_en(rlydiag4_oc_rly9_en),
    .rlydiag4_oc_rly9_in(rlydiag4_oc_rly9_in),
    // RlyDiag4.SCG_VLV1
    .rlydiag4_scg_vlv1_en(rlydiag4_scg_vlv1_en),
    .rlydiag4_scg_vlv1_in(rlydiag4_scg_vlv1_in),
    // RlyDiag4.OL_VLV1
    .rlydiag4_ol_vlv1_en(rlydiag4_ol_vlv1_en),
    .rlydiag4_ol_vlv1_in(rlydiag4_ol_vlv1_in),
    // RlyDiag4.TSD_VLV1
    .rlydiag4_tsd_vlv1_en(rlydiag4_tsd_vlv1_en),
    .rlydiag4_tsd_vlv1_in(rlydiag4_tsd_vlv1_in),
    // RlyDiag4.OC_VLV1
    .rlydiag4_oc_vlv1_en(rlydiag4_oc_vlv1_en),
    .rlydiag4_oc_vlv1_in(rlydiag4_oc_vlv1_in),

    // VlvDiag.SCG_VLV2
    .vlvdiag_scg_vlv2_en(vlvdiag_scg_vlv2_en),
    .vlvdiag_scg_vlv2_in(vlvdiag_scg_vlv2_in),
    // VlvDiag.OL_VLV2
    .vlvdiag_ol_vlv2_en(vlvdiag_ol_vlv2_en),
    .vlvdiag_ol_vlv2_in(vlvdiag_ol_vlv2_in),
    // VlvDiag.TSD_VLV2
    .vlvdiag_tsd_vlv2_en(vlvdiag_tsd_vlv2_en),
    .vlvdiag_tsd_vlv2_in(vlvdiag_tsd_vlv2_in),
    // VlvDiag.OC_VLV2
    .vlvdiag_oc_vlv2_en(vlvdiag_oc_vlv2_en),
    .vlvdiag_oc_vlv2_in(vlvdiag_oc_vlv2_in),
    // VlvDiag.SCG_VLV3
    .vlvdiag_scg_vlv3_en(vlvdiag_scg_vlv3_en),
    .vlvdiag_scg_vlv3_in(vlvdiag_scg_vlv3_in),
    // VlvDiag.OL_VLV3
    .vlvdiag_ol_vlv3_en(vlvdiag_ol_vlv3_en),
    .vlvdiag_ol_vlv3_in(vlvdiag_ol_vlv3_in),
    // VlvDiag.TSD_VLV3
    .vlvdiag_tsd_vlv3_en(vlvdiag_tsd_vlv3_en),
    .vlvdiag_tsd_vlv3_in(vlvdiag_tsd_vlv3_in),
    // VlvDiag.OC_VLV3
    .vlvdiag_oc_vlv3_en(vlvdiag_oc_vlv3_en),
    .vlvdiag_oc_vlv3_in(vlvdiag_oc_vlv3_in),

    // HbDiag0.TSD_HS1
    .hbdiag0_tsd_hs1_en(hbdiag0_tsd_hs1_en),
    .hbdiag0_tsd_hs1_in(hbdiag0_tsd_hs1_in),
    // HbDiag0.OC_HS1
    .hbdiag0_oc_hs1_en(hbdiag0_oc_hs1_en),
    .hbdiag0_oc_hs1_in(hbdiag0_oc_hs1_in),
    // HbDiag0.TSD_LS1
    .hbdiag0_tsd_ls1_en(hbdiag0_tsd_ls1_en),
    .hbdiag0_tsd_ls1_in(hbdiag0_tsd_ls1_in),
    // HbDiag0.OC_LS1
    .hbdiag0_oc_ls1_en(hbdiag0_oc_ls1_en),
    .hbdiag0_oc_ls1_in(hbdiag0_oc_ls1_in),
    // HbDiag0.SCG_HB1
    .hbdiag0_scg_hb1_en(hbdiag0_scg_hb1_en),
    .hbdiag0_scg_hb1_in(hbdiag0_scg_hb1_in),
    // HbDiag0.SCB_HB1
    .hbdiag0_scb_hb1_en(hbdiag0_scb_hb1_en),
    .hbdiag0_scb_hb1_in(hbdiag0_scb_hb1_in),
    // HbDiag0.OL_HB1
    .hbdiag0_ol_hb1_en(hbdiag0_ol_hb1_en),
    .hbdiag0_ol_hb1_in(hbdiag0_ol_hb1_in),

    // HbDiag1.TSD_HS2
    .hbdiag1_tsd_hs2_en(hbdiag1_tsd_hs2_en),
    .hbdiag1_tsd_hs2_in(hbdiag1_tsd_hs2_in),
    // HbDiag1.OC_HS2
    .hbdiag1_oc_hs2_en(hbdiag1_oc_hs2_en),
    .hbdiag1_oc_hs2_in(hbdiag1_oc_hs2_in),
    // HbDiag1.TSD_LS2
    .hbdiag1_tsd_ls2_en(hbdiag1_tsd_ls2_en),
    .hbdiag1_tsd_ls2_in(hbdiag1_tsd_ls2_in),
    // HbDiag1.OC_LS2
    .hbdiag1_oc_ls2_en(hbdiag1_oc_ls2_en),
    .hbdiag1_oc_ls2_in(hbdiag1_oc_ls2_in),
    // HbDiag1.SCG_HB2
    .hbdiag1_scg_hb2_en(hbdiag1_scg_hb2_en),
    .hbdiag1_scg_hb2_in(hbdiag1_scg_hb2_in),
    // HbDiag1.SCB_HB2
    .hbdiag1_scb_hb2_en(hbdiag1_scb_hb2_en),
    .hbdiag1_scb_hb2_in(hbdiag1_scb_hb2_in),
    // HbDiag1.OL_HB2
    .hbdiag1_ol_hb2_en(hbdiag1_ol_hb2_en),
    .hbdiag1_ol_hb2_in(hbdiag1_ol_hb2_in),

    // RstDiag.RSTB_EVENT
    .rstdiag_rstb_event_en(rstdiag_rstb_event_en),
    .rstdiag_rstb_event_in(rstdiag_rstb_event_in),
    // RstDiag.WD_RST_EVENT
    .rstdiag_wd_rst_event_en(rstdiag_wd_rst_event_en),
    .rstdiag_wd_rst_event_in(rstdiag_wd_rst_event_in),
    // RstDiag.SOFTWARE_RST_EVENT
    .rstdiag_software_rst_event_en(rstdiag_software_rst_event_en),
    .rstdiag_software_rst_event_in(rstdiag_software_rst_event_in),
    // RstDiag.VDD5_UV_RST_EVENT
    .rstdiag_vdd5_uv_rst_event_en(rstdiag_vdd5_uv_rst_event_en),
    .rstdiag_vdd5_uv_rst_event_in(rstdiag_vdd5_uv_rst_event_in),
    // RstDiag.VDD5_OV_RST_EVENT
    .rstdiag_vdd5_ov_rst_event_en(rstdiag_vdd5_ov_rst_event_en),
    .rstdiag_vdd5_ov_rst_event_in(rstdiag_vdd5_ov_rst_event_in),
    // RstDiag.POR_EVENT
    .rstdiag_por_event_en(rstdiag_por_event_en),
    .rstdiag_por_event_in(rstdiag_por_event_in),

    // GLBStatus.TSD_OC_FAIL
    .glbstatus_tsd_oc_fail_en(glbstatus_tsd_oc_fail_en),
    .glbstatus_tsd_oc_fail_in(glbstatus_tsd_oc_fail_in),
    // GLBStatus.SC_OL_FAIL
    .glbstatus_sc_ol_fail_en(glbstatus_sc_ol_fail_en),
    .glbstatus_sc_ol_fail_in(glbstatus_sc_ol_fail_in),
    // GLBStatus.WD_SV_FAIL
    .glbstatus_wd_sv_fail_en(glbstatus_wd_sv_fail_en),
    .glbstatus_wd_sv_fail_in(glbstatus_wd_sv_fail_in),
    // GLBStatus.SUP_FAIL_DIS_DRV
    .glbstatus_sup_fail_dis_drv_en(glbstatus_sup_fail_dis_drv_en),
    .glbstatus_sup_fail_dis_drv_in(glbstatus_sup_fail_dis_drv_in),
    // GLBStatus.VRS_FAIL
    .glbstatus_vrs_fail_en(glbstatus_vrs_fail_en),
    .glbstatus_vrs_fail_in(glbstatus_vrs_fail_in),
    // GLBStatus.OTP_FAIL
    .glbstatus_otp_fail_en(glbstatus_otp_fail_en),
    .glbstatus_otp_fail_in(glbstatus_otp_fail_in),
    // GLBStatus.SPI_MSC_FAIL
    .glbstatus_spi_msc_fail_en(glbstatus_spi_msc_fail_en),
    .glbstatus_spi_msc_fail_in(glbstatus_spi_msc_fail_in),
    // GLBStatus.GND_FAIL
    .glbstatus_gnd_fail_en(glbstatus_gnd_fail_en),
    .glbstatus_gnd_fail_in(glbstatus_gnd_fail_in),

    // WdQuestion.LFSR
    .wdquestion_lfsr_en(wdquestion_lfsr_en),
    .wdquestion_lfsr_in(wdquestion_lfsr_in),

    // WdPassCnt.WD_RFH_CNT
    .wdpasscnt_wd_rfh_cnt_en(wdpasscnt_wd_rfh_cnt_en),
    .wdpasscnt_wd_rfh_cnt_in(wdpasscnt_wd_rfh_cnt_in),

    // WdFailCnt.WD_ERR_CNT
    .wdfailcnt_wd_err_cnt_en(wdfailcnt_wd_err_cnt_en),
    .wdfailcnt_wd_err_cnt_in(wdfailcnt_wd_err_cnt_in),
    // WdFailCnt.RST_ERR_CNT
    .wdfailcnt_rst_err_cnt_en(wdfailcnt_rst_err_cnt_en),
    .wdfailcnt_rst_err_cnt_in(wdfailcnt_rst_err_cnt_in),

    // PSState0.OUT_STATE_IGN
    .psstate0_out_state_ign_en(psstate0_out_state_ign_en),
    .psstate0_out_state_ign_in(psstate0_out_state_ign_in),
    // PSState0.OUT_STATE_INJ
    .psstate0_out_state_inj_en(psstate0_out_state_inj_en),
    .psstate0_out_state_inj_in(psstate0_out_state_inj_in),

    // PSState1.OUT_STATE_RLY
    .psstate1_out_state_rly_en(psstate1_out_state_rly_en),
    .psstate1_out_state_rly_in(psstate1_out_state_rly_in),

    // PSState2.OUT_STATE_RLY
    .psstate2_out_state_rly_en(psstate2_out_state_rly_en),
    .psstate2_out_state_rly_in(psstate2_out_state_rly_in),
    // PSState2.OUT_STATE_HTR
    .psstate2_out_state_htr_en(psstate2_out_state_htr_en),
    .psstate2_out_state_htr_in(psstate2_out_state_htr_in),
    // PSState2.OUT_STATE_VLV
    .psstate2_out_state_vlv_en(psstate2_out_state_vlv_en),
    .psstate2_out_state_vlv_in(psstate2_out_state_vlv_in),

    // PSState3.OUT_STATE_HS
    .psstate3_out_state_hs_en(psstate3_out_state_hs_en),
    .psstate3_out_state_hs_in(psstate3_out_state_hs_in),
    // PSState3.OUT_STATE_LS
    .psstate3_out_state_ls_en(psstate3_out_state_ls_en),
    .psstate3_out_state_ls_in(psstate3_out_state_ls_in),

    // InState0.DIN
    .instate0_din_en(instate0_din_en),
    .instate0_din_in(instate0_din_in),

    // InState1.DIN
    .instate1_din_en(instate1_din_en),
    .instate1_din_in(instate1_din_in),

    // EnState0.OE
    .enstate0_oe_en(enstate0_oe_en),
    .enstate0_oe_in(enstate0_oe_in),
    // EnState0.DEN_RLY
    .enstate0_den_rly_en(enstate0_den_rly_en),
    .enstate0_den_rly_in(enstate0_den_rly_in),
    // EnState0.DEN_DRV
    .enstate0_den_drv_en(enstate0_den_drv_en),
    .enstate0_den_drv_in(enstate0_den_drv_in),
    // EnState0.DNDIS_DRV
    .enstate0_dndis_drv_en(enstate0_dndis_drv_en),
    .enstate0_dndis_drv_in(enstate0_dndis_drv_in),

    // MaskID.MASK_ID
    .maskid_mask_id_en(maskid_mask_id_en),
    .maskid_mask_id_in(maskid_mask_id_in),

    // Cmd0.Code
    .cmd0_code_out(cmd0_code_out),

    // CmdWdCheck.MCU_REPLY
    .cmdwdcheck_mcu_reply_out(cmdwdcheck_mcu_reply_out),

    // CmdWdLdSd.SEED
    .cmdwdldsd_seed_out(cmdwdldsd_seed_out),

    // CmdSoftRst.SOFTWARE_RST
    .cmdsoftrst_software_rst_out(cmdsoftrst_software_rst_out),

    // MscRCmd0.DisDrvConfig0
    .mscrcmd0_disdrvconfig0_out(mscrcmd0_disdrvconfig0_out),
    // MscRCmd0.DisDrvConfig1
    .mscrcmd0_disdrvconfig1_out(mscrcmd0_disdrvconfig1_out),
    // MscRCmd0.DisDrvConfig2
    .mscrcmd0_disdrvconfig2_out(mscrcmd0_disdrvconfig2_out),
    // MscRCmd0.DenConfig0
    .mscrcmd0_denconfig0_out(mscrcmd0_denconfig0_out),
    // MscRCmd0.DenConfig1
    .mscrcmd0_denconfig1_out(mscrcmd0_denconfig1_out),
    // MscRCmd0.DenConfig2
    .mscrcmd0_denconfig2_out(mscrcmd0_denconfig2_out),
    // MscRCmd0.DenConfig3
    .mscrcmd0_denconfig3_out(mscrcmd0_denconfig3_out),
    // MscRCmd0.DenConfig4
    .mscrcmd0_denconfig4_out(mscrcmd0_denconfig4_out),

    // MscRCmd1.OEConfig0
    .mscrcmd1_oeconfig0_out(mscrcmd1_oeconfig0_out),
    // MscRCmd1.OEConfig1
    .mscrcmd1_oeconfig1_out(mscrcmd1_oeconfig1_out),
    // MscRCmd1.OEConfig2
    .mscrcmd1_oeconfig2_out(mscrcmd1_oeconfig2_out),
    // MscRCmd1.OEConfig3
    .mscrcmd1_oeconfig3_out(mscrcmd1_oeconfig3_out),
    // MscRCmd1.Cont0
    .mscrcmd1_cont0_out(mscrcmd1_cont0_out),
    // MscRCmd1.Cont1
    .mscrcmd1_cont1_out(mscrcmd1_cont1_out),
    // MscRCmd1.Cont2
    .mscrcmd1_cont2_out(mscrcmd1_cont2_out),

    // MscRCmd2.DDConfig0
    .mscrcmd2_ddconfig0_out(mscrcmd2_ddconfig0_out),
    // MscRCmd2.DDConfig1
    .mscrcmd2_ddconfig1_out(mscrcmd2_ddconfig1_out),
    // MscRCmd2.DDConfig2
    .mscrcmd2_ddconfig2_out(mscrcmd2_ddconfig2_out),
    // MscRCmd2.BRIConfig
    .mscrcmd2_briconfig_out(mscrcmd2_briconfig_out),
    // MscRCmd2.DlyOffConfig
    .mscrcmd2_dlyoffconfig_out(mscrcmd2_dlyoffconfig_out),
    // MscRCmd2.CurrLimConfig0
    .mscrcmd2_currlimconfig0_out(mscrcmd2_currlimconfig0_out),
    // MscRCmd2.CurrLimConfig1
    .mscrcmd2_currlimconfig1_out(mscrcmd2_currlimconfig1_out),
    // MscRCmd2.CurrLimConfig2
    .mscrcmd2_currlimconfig2_out(mscrcmd2_currlimconfig2_out),

    // MscRCmd3.OutDiagConfig0
    .mscrcmd3_outdiagconfig0_out(mscrcmd3_outdiagconfig0_out),
    // MscRCmd3.OutDiagConfig1
    .mscrcmd3_outdiagconfig1_out(mscrcmd3_outdiagconfig1_out),
    // MscRCmd3.OutDiagConfig2
    .mscrcmd3_outdiagconfig2_out(mscrcmd3_outdiagconfig2_out),
    // MscRCmd3.OutDiagConfig3
    .mscrcmd3_outdiagconfig3_out(mscrcmd3_outdiagconfig3_out),
    // MscRCmd3.OutDiagConfig4
    .mscrcmd3_outdiagconfig4_out(mscrcmd3_outdiagconfig4_out),
    // MscRCmd3.IgnDiagConfig
    .mscrcmd3_igndiagconfig_out(mscrcmd3_igndiagconfig_out),

    // MscRCmd4.DinConfig0
    .mscrcmd4_dinconfig0_out(mscrcmd4_dinconfig0_out),
    // MscRCmd4.DinConfig1
    .mscrcmd4_dinconfig1_out(mscrcmd4_dinconfig1_out),
    // MscRCmd4.DinConfig2
    .mscrcmd4_dinconfig2_out(mscrcmd4_dinconfig2_out),
    // MscRCmd4.DinConfig3
    .mscrcmd4_dinconfig3_out(mscrcmd4_dinconfig3_out),
    // MscRCmd4.DinConfig4
    .mscrcmd4_dinconfig4_out(mscrcmd4_dinconfig4_out),
    // MscRCmd4.DinConfig5
    .mscrcmd4_dinconfig5_out(mscrcmd4_dinconfig5_out),
    // MscRCmd4.DinConfig6
    .mscrcmd4_dinconfig6_out(mscrcmd4_dinconfig6_out),
    // MscRCmd4.DinConfig7
    .mscrcmd4_dinconfig7_out(mscrcmd4_dinconfig7_out),

    // MscRCmd5.DinConfig8
    .mscrcmd5_dinconfig8_out(mscrcmd5_dinconfig8_out),
    // MscRCmd5.DinConfig9
    .mscrcmd5_dinconfig9_out(mscrcmd5_dinconfig9_out),
    // MscRCmd5.DinConfig10
    .mscrcmd5_dinconfig10_out(mscrcmd5_dinconfig10_out),
    // MscRCmd5.DinConfig11
    .mscrcmd5_dinconfig11_out(mscrcmd5_dinconfig11_out),
    // MscRCmd5.RstbConfig
    .mscrcmd5_rstbconfig_out(mscrcmd5_rstbconfig_out),
    // MscRCmd5.FaultbConfig0
    .mscrcmd5_faultbconfig0_out(mscrcmd5_faultbconfig0_out),
    // MscRCmd5.FaultbConfig1
    .mscrcmd5_faultbconfig1_out(mscrcmd5_faultbconfig1_out),
    // MscRCmd5.FaultbConfig2
    .mscrcmd5_faultbconfig2_out(mscrcmd5_faultbconfig2_out),

    // MscRCmd6.WDConfig0
    .mscrcmd6_wdconfig0_out(mscrcmd6_wdconfig0_out),
    // MscRCmd6.WDConfig1
    .mscrcmd6_wdconfig1_out(mscrcmd6_wdconfig1_out),
    // MscRCmd6.VrsConfig0
    .mscrcmd6_vrsconfig0_out(mscrcmd6_vrsconfig0_out),
    // MscRCmd6.VrsConfig1
    .mscrcmd6_vrsconfig1_out(mscrcmd6_vrsconfig1_out),
    // MscRCmd6.VrsConfig2
    .mscrcmd6_vrsconfig2_out(mscrcmd6_vrsconfig2_out),
    // MscRCmd6.MscConfig0
    .mscrcmd6_mscconfig0_out(mscrcmd6_mscconfig0_out),
    // MscRCmd6.MscConfig1
    .mscrcmd6_mscconfig1_out(mscrcmd6_mscconfig1_out),
    // MscRCmd6.AoutConfig
    .mscrcmd6_aoutconfig_out(mscrcmd6_aoutconfig_out),

    // MscRCmd7.VrsDiag
    .mscrcmd7_vrsdiag_out(mscrcmd7_vrsdiag_out),
    // MscRCmd7.SupDiag
    .mscrcmd7_supdiag_out(mscrcmd7_supdiag_out),
    // MscRCmd7.ExtDiag0
    .mscrcmd7_extdiag0_out(mscrcmd7_extdiag0_out),
    // MscRCmd7.ExtDiag1
    .mscrcmd7_extdiag1_out(mscrcmd7_extdiag1_out),

    // MscRCmd8.InjDiag0
    .mscrcmd8_injdiag0_out(mscrcmd8_injdiag0_out),
    // MscRCmd8.InjDiag1
    .mscrcmd8_injdiag1_out(mscrcmd8_injdiag1_out),
    // MscRCmd8.IgnDiag0
    .mscrcmd8_igndiag0_out(mscrcmd8_igndiag0_out),
    // MscRCmd8.IgnDiag1
    .mscrcmd8_igndiag1_out(mscrcmd8_igndiag1_out),
    // MscRCmd8.HbDiag0
    .mscrcmd8_hbdiag0_out(mscrcmd8_hbdiag0_out),
    // MscRCmd8.HbDiag1
    .mscrcmd8_hbdiag1_out(mscrcmd8_hbdiag1_out),

    // MscRCmd9.RlyDiag0
    .mscrcmd9_rlydiag0_out(mscrcmd9_rlydiag0_out),
    // MscRCmd9.RlyDiag1
    .mscrcmd9_rlydiag1_out(mscrcmd9_rlydiag1_out),
    // MscRCmd9.RlyDiag2
    .mscrcmd9_rlydiag2_out(mscrcmd9_rlydiag2_out),
    // MscRCmd9.RlyDiag3
    .mscrcmd9_rlydiag3_out(mscrcmd9_rlydiag3_out),
    // MscRCmd9.RlyDiag4
    .mscrcmd9_rlydiag4_out(mscrcmd9_rlydiag4_out),
    // MscRCmd9.HtrDiag0
    .mscrcmd9_htrdiag0_out(mscrcmd9_htrdiag0_out),
    // MscRCmd9.VlvDiag
    .mscrcmd9_vlvdiag_out(mscrcmd9_vlvdiag_out),
    // MscRCmd9.RstDiag
    .mscrcmd9_rstdiag_out(mscrcmd9_rstdiag_out),

    // MscRCmd10.GLBStatus
    .mscrcmd10_glbstatus_out(mscrcmd10_glbstatus_out),
    // MscRCmd10.WdQuestion
    .mscrcmd10_wdquestion_out(mscrcmd10_wdquestion_out),
    // MscRCmd10.WdPassCnt
    .mscrcmd10_wdpasscnt_out(mscrcmd10_wdpasscnt_out),
    // MscRCmd10.WdFailCnt
    .mscrcmd10_wdfailcnt_out(mscrcmd10_wdfailcnt_out),

    // MscRCmd11.PSState0
    .mscrcmd11_psstate0_out(mscrcmd11_psstate0_out),
    // MscRCmd11.PSState1
    .mscrcmd11_psstate1_out(mscrcmd11_psstate1_out),
    // MscRCmd11.PSState2
    .mscrcmd11_psstate2_out(mscrcmd11_psstate2_out),
    // MscRCmd11.PSState3
    .mscrcmd11_psstate3_out(mscrcmd11_psstate3_out),
    // MscRCmd11.InState0
    .mscrcmd11_instate0_out(mscrcmd11_instate0_out),
    // MscRCmd11.InState1
    .mscrcmd11_instate1_out(mscrcmd11_instate1_out),
    // MscRCmd11.EnState0
    .mscrcmd11_enstate0_out(mscrcmd11_enstate0_out),
    // MscRCmd11.MaskId
    .mscrcmd11_maskid_out(mscrcmd11_maskid_out),

    // CmdSpecialMode.SM_DIS_TSD
    .cmdspecialmode_sm_dis_tsd_en(cmdspecialmode_sm_dis_tsd_en),
    .cmdspecialmode_sm_dis_tsd_in(cmdspecialmode_sm_dis_tsd_in),
    .cmdspecialmode_sm_dis_tsd_out(cmdspecialmode_sm_dis_tsd_out),
    // CmdSpecialMode.SM_DIS_VDD5_UV
    .cmdspecialmode_sm_dis_vdd5_uv_en(cmdspecialmode_sm_dis_vdd5_uv_en),
    .cmdspecialmode_sm_dis_vdd5_uv_in(cmdspecialmode_sm_dis_vdd5_uv_in),
    .cmdspecialmode_sm_dis_vdd5_uv_out(cmdspecialmode_sm_dis_vdd5_uv_out),
    // CmdSpecialMode.SM_DIS_VDD5_OV
    .cmdspecialmode_sm_dis_vdd5_ov_en(cmdspecialmode_sm_dis_vdd5_ov_en),
    .cmdspecialmode_sm_dis_vdd5_ov_in(cmdspecialmode_sm_dis_vdd5_ov_in),
    .cmdspecialmode_sm_dis_vdd5_ov_out(cmdspecialmode_sm_dis_vdd5_ov_out),
    // CmdSpecialMode.SM_DIS_VPWR_OV
    .cmdspecialmode_sm_dis_vpwr_ov_en(cmdspecialmode_sm_dis_vpwr_ov_en),
    .cmdspecialmode_sm_dis_vpwr_ov_in(cmdspecialmode_sm_dis_vpwr_ov_in),
    .cmdspecialmode_sm_dis_vpwr_ov_out(cmdspecialmode_sm_dis_vpwr_ov_out),
    // CmdSpecialMode.SM_DIS_VPWR_UV
    .cmdspecialmode_sm_dis_vpwr_uv_en(cmdspecialmode_sm_dis_vpwr_uv_en),
    .cmdspecialmode_sm_dis_vpwr_uv_in(cmdspecialmode_sm_dis_vpwr_uv_in),
    .cmdspecialmode_sm_dis_vpwr_uv_out(cmdspecialmode_sm_dis_vpwr_uv_out),
    // CmdSpecialMode.SM_DIS_VCP_UV
    .cmdspecialmode_sm_dis_vcp_uv_en(cmdspecialmode_sm_dis_vcp_uv_en),
    .cmdspecialmode_sm_dis_vcp_uv_in(cmdspecialmode_sm_dis_vcp_uv_in),
    .cmdspecialmode_sm_dis_vcp_uv_out(cmdspecialmode_sm_dis_vcp_uv_out),
    // CmdSpecialMode.SM_DIS_OC
    .cmdspecialmode_sm_dis_oc_en(cmdspecialmode_sm_dis_oc_en),
    .cmdspecialmode_sm_dis_oc_in(cmdspecialmode_sm_dis_oc_in),
    .cmdspecialmode_sm_dis_oc_out(cmdspecialmode_sm_dis_oc_out),
    // CmdSpecialMode.SM_DIS_IGN_SCG_GNDLOSS
    .cmdspecialmode_sm_dis_ign_scg_gndloss_en(cmdspecialmode_sm_dis_ign_scg_gndloss_en),
    .cmdspecialmode_sm_dis_ign_scg_gndloss_in(cmdspecialmode_sm_dis_ign_scg_gndloss_in),
    .cmdspecialmode_sm_dis_ign_scg_gndloss_out(cmdspecialmode_sm_dis_ign_scg_gndloss_out),

    // CmdTM.TM_CODE
    .cmdtm_tm_code_en(cmdtm_tm_code_en),
    .cmdtm_tm_code_in(cmdtm_tm_code_in),
    .cmdtm_tm_code_out(cmdtm_tm_code_out),

    // PageVrb.CODE
    .pagevrb_code_en(pagevrb_code_en),
    .pagevrb_code_in(pagevrb_code_in),
    .pagevrb_code_out(pagevrb_code_out),

    // Local Bus
    .waddr(waddr),
    .wdata(wdata),
    .wen(wen),
    .wstrb(wstrb),
    .wready(wready),
    .raddr(raddr),
    .ren(ren),
    .rdata(rdata),
    .rvalid(rvalid)
    );