// Created with regmapGen v1.0.3

package Uchip_regmap0_pkg;

parameter BASE_ADDR = 0;
parameter DATA_WIDTH = 8;
parameter ADDR_WIDTH = 8;

// DisDrvConfig0
parameter DISDRVCONFIG0_ADDR = 8'h0;
parameter DISDRVCONFIG0_RESET = 8'hff;

// DisDrvConfig0.DDIS_DRVB_CFG_INJ
parameter DISDRVCONFIG0_DDIS_DRVB_CFG_INJ_WIDTH = 4;
parameter DISDRVCONFIG0_DDIS_DRVB_CFG_INJ_LSB = 0;
parameter DISDRVCONFIG0_DDIS_DRVB_CFG_INJ_MASK = 8'hf;
parameter DISDRVCONFIG0_DDIS_DRVB_CFG_INJ_RESET = 4'hf;

// DisDrvConfig0.DDIS_DRVB_CFG_IGN
parameter DISDRVCONFIG0_DDIS_DRVB_CFG_IGN_WIDTH = 4;
parameter DISDRVCONFIG0_DDIS_DRVB_CFG_IGN_LSB = 4;
parameter DISDRVCONFIG0_DDIS_DRVB_CFG_IGN_MASK = 8'hf0;
parameter DISDRVCONFIG0_DDIS_DRVB_CFG_IGN_RESET = 4'hf;


// DisDrvConfig1
parameter DISDRVCONFIG1_ADDR = 8'h1;
parameter DISDRVCONFIG1_RESET = 8'hff;

// DisDrvConfig1.DDIS_DRVB_CFG_RLY
parameter DISDRVCONFIG1_DDIS_DRVB_CFG_RLY_WIDTH = 8;
parameter DISDRVCONFIG1_DDIS_DRVB_CFG_RLY_LSB = 0;
parameter DISDRVCONFIG1_DDIS_DRVB_CFG_RLY_MASK = 8'hff;
parameter DISDRVCONFIG1_DDIS_DRVB_CFG_RLY_RESET = 8'hff;


// DisDrvConfig2
parameter DISDRVCONFIG2_ADDR = 8'h2;
parameter DISDRVCONFIG2_RESET = 8'hff;

// DisDrvConfig2.DDIS_DRVB_CFG_RLY
parameter DISDRVCONFIG2_DDIS_DRVB_CFG_RLY_WIDTH = 1;
parameter DISDRVCONFIG2_DDIS_DRVB_CFG_RLY_LSB = 0;
parameter DISDRVCONFIG2_DDIS_DRVB_CFG_RLY_MASK = 8'h1;
parameter DISDRVCONFIG2_DDIS_DRVB_CFG_RLY_RESET = 1'h1;

// DisDrvConfig2.DDIS_DRVB_CFG_VLV
parameter DISDRVCONFIG2_DDIS_DRVB_CFG_VLV_WIDTH = 3;
parameter DISDRVCONFIG2_DDIS_DRVB_CFG_VLV_LSB = 1;
parameter DISDRVCONFIG2_DDIS_DRVB_CFG_VLV_MASK = 8'he;
parameter DISDRVCONFIG2_DDIS_DRVB_CFG_VLV_RESET = 3'h7;

// DisDrvConfig2.DDIS_DRVB_CFG_HTR
parameter DISDRVCONFIG2_DDIS_DRVB_CFG_HTR_WIDTH = 2;
parameter DISDRVCONFIG2_DDIS_DRVB_CFG_HTR_LSB = 4;
parameter DISDRVCONFIG2_DDIS_DRVB_CFG_HTR_MASK = 8'h30;
parameter DISDRVCONFIG2_DDIS_DRVB_CFG_HTR_RESET = 2'h3;

// DisDrvConfig2.DDIS_DRVB_CFG_HB
parameter DISDRVCONFIG2_DDIS_DRVB_CFG_HB_WIDTH = 2;
parameter DISDRVCONFIG2_DDIS_DRVB_CFG_HB_LSB = 6;
parameter DISDRVCONFIG2_DDIS_DRVB_CFG_HB_MASK = 8'hc0;
parameter DISDRVCONFIG2_DDIS_DRVB_CFG_HB_RESET = 2'h3;


// DenConfig0
parameter DENCONFIG0_ADDR = 8'h3;
parameter DENCONFIG0_RESET = 8'hf;

// DenConfig0.DEN_DRV_CFG_IGN
parameter DENCONFIG0_DEN_DRV_CFG_IGN_WIDTH = 4;
parameter DENCONFIG0_DEN_DRV_CFG_IGN_LSB = 0;
parameter DENCONFIG0_DEN_DRV_CFG_IGN_MASK = 8'hf;
parameter DENCONFIG0_DEN_DRV_CFG_IGN_RESET = 4'hf;


// DenConfig1
parameter DENCONFIG1_ADDR = 8'h4;
parameter DENCONFIG1_RESET = 8'h1f;

// DenConfig1.DEN_DRV_CFG_RLY1
parameter DENCONFIG1_DEN_DRV_CFG_RLY1_WIDTH = 1;
parameter DENCONFIG1_DEN_DRV_CFG_RLY1_LSB = 0;
parameter DENCONFIG1_DEN_DRV_CFG_RLY1_MASK = 8'h1;
parameter DENCONFIG1_DEN_DRV_CFG_RLY1_RESET = 1'h1;

// DenConfig1.DEN_RLY_CFG_RLY1
parameter DENCONFIG1_DEN_RLY_CFG_RLY1_WIDTH = 1;
parameter DENCONFIG1_DEN_RLY_CFG_RLY1_LSB = 1;
parameter DENCONFIG1_DEN_RLY_CFG_RLY1_MASK = 8'h2;
parameter DENCONFIG1_DEN_RLY_CFG_RLY1_RESET = 1'h1;

// DenConfig1.DEN_DRV_CFG_RLY2
parameter DENCONFIG1_DEN_DRV_CFG_RLY2_WIDTH = 1;
parameter DENCONFIG1_DEN_DRV_CFG_RLY2_LSB = 2;
parameter DENCONFIG1_DEN_DRV_CFG_RLY2_MASK = 8'h4;
parameter DENCONFIG1_DEN_DRV_CFG_RLY2_RESET = 1'h1;

// DenConfig1.DEN_RLY_CFG_RLY2
parameter DENCONFIG1_DEN_RLY_CFG_RLY2_WIDTH = 1;
parameter DENCONFIG1_DEN_RLY_CFG_RLY2_LSB = 3;
parameter DENCONFIG1_DEN_RLY_CFG_RLY2_MASK = 8'h8;
parameter DENCONFIG1_DEN_RLY_CFG_RLY2_RESET = 1'h1;

// DenConfig1.DEN_DRV_CFG_RLY3
parameter DENCONFIG1_DEN_DRV_CFG_RLY3_WIDTH = 1;
parameter DENCONFIG1_DEN_DRV_CFG_RLY3_LSB = 4;
parameter DENCONFIG1_DEN_DRV_CFG_RLY3_MASK = 8'h10;
parameter DENCONFIG1_DEN_DRV_CFG_RLY3_RESET = 1'h1;

// DenConfig1.DEN_RLY_CFG_RLY3
parameter DENCONFIG1_DEN_RLY_CFG_RLY3_WIDTH = 1;
parameter DENCONFIG1_DEN_RLY_CFG_RLY3_LSB = 5;
parameter DENCONFIG1_DEN_RLY_CFG_RLY3_MASK = 8'h20;
parameter DENCONFIG1_DEN_RLY_CFG_RLY3_RESET = 1'h0;

// DenConfig1.DEN_DRV_CFG_RLY4
parameter DENCONFIG1_DEN_DRV_CFG_RLY4_WIDTH = 1;
parameter DENCONFIG1_DEN_DRV_CFG_RLY4_LSB = 6;
parameter DENCONFIG1_DEN_DRV_CFG_RLY4_MASK = 8'h40;
parameter DENCONFIG1_DEN_DRV_CFG_RLY4_RESET = 1'h0;

// DenConfig1.DEN_RLY_CFG_RLY4
parameter DENCONFIG1_DEN_RLY_CFG_RLY4_WIDTH = 1;
parameter DENCONFIG1_DEN_RLY_CFG_RLY4_LSB = 7;
parameter DENCONFIG1_DEN_RLY_CFG_RLY4_MASK = 8'h80;
parameter DENCONFIG1_DEN_RLY_CFG_RLY4_RESET = 1'h0;


// DenConfig2
parameter DENCONFIG2_ADDR = 8'h5;
parameter DENCONFIG2_RESET = 8'h0;

// DenConfig2.DEN_DRV_CFG_RLY5
parameter DENCONFIG2_DEN_DRV_CFG_RLY5_WIDTH = 1;
parameter DENCONFIG2_DEN_DRV_CFG_RLY5_LSB = 0;
parameter DENCONFIG2_DEN_DRV_CFG_RLY5_MASK = 8'h1;
parameter DENCONFIG2_DEN_DRV_CFG_RLY5_RESET = 1'h0;

// DenConfig2.DEN_RLY_CFG_RLY5
parameter DENCONFIG2_DEN_RLY_CFG_RLY5_WIDTH = 1;
parameter DENCONFIG2_DEN_RLY_CFG_RLY5_LSB = 1;
parameter DENCONFIG2_DEN_RLY_CFG_RLY5_MASK = 8'h2;
parameter DENCONFIG2_DEN_RLY_CFG_RLY5_RESET = 1'h0;

// DenConfig2.DEN_DRV_CFG_RLY6
parameter DENCONFIG2_DEN_DRV_CFG_RLY6_WIDTH = 1;
parameter DENCONFIG2_DEN_DRV_CFG_RLY6_LSB = 2;
parameter DENCONFIG2_DEN_DRV_CFG_RLY6_MASK = 8'h4;
parameter DENCONFIG2_DEN_DRV_CFG_RLY6_RESET = 1'h0;

// DenConfig2.DEN_RLY_CFG_RLY6
parameter DENCONFIG2_DEN_RLY_CFG_RLY6_WIDTH = 1;
parameter DENCONFIG2_DEN_RLY_CFG_RLY6_LSB = 3;
parameter DENCONFIG2_DEN_RLY_CFG_RLY6_MASK = 8'h8;
parameter DENCONFIG2_DEN_RLY_CFG_RLY6_RESET = 1'h0;

// DenConfig2.DEN_DRV_CFG_RLY7
parameter DENCONFIG2_DEN_DRV_CFG_RLY7_WIDTH = 1;
parameter DENCONFIG2_DEN_DRV_CFG_RLY7_LSB = 4;
parameter DENCONFIG2_DEN_DRV_CFG_RLY7_MASK = 8'h10;
parameter DENCONFIG2_DEN_DRV_CFG_RLY7_RESET = 1'h0;

// DenConfig2.DEN_RLY_CFG_RLY7
parameter DENCONFIG2_DEN_RLY_CFG_RLY7_WIDTH = 1;
parameter DENCONFIG2_DEN_RLY_CFG_RLY7_LSB = 5;
parameter DENCONFIG2_DEN_RLY_CFG_RLY7_MASK = 8'h20;
parameter DENCONFIG2_DEN_RLY_CFG_RLY7_RESET = 1'h0;

// DenConfig2.DEN_DRV_CFG_RLY8
parameter DENCONFIG2_DEN_DRV_CFG_RLY8_WIDTH = 1;
parameter DENCONFIG2_DEN_DRV_CFG_RLY8_LSB = 6;
parameter DENCONFIG2_DEN_DRV_CFG_RLY8_MASK = 8'h40;
parameter DENCONFIG2_DEN_DRV_CFG_RLY8_RESET = 1'h0;

// DenConfig2.DEN_RLY_CFG_RLY8
parameter DENCONFIG2_DEN_RLY_CFG_RLY8_WIDTH = 1;
parameter DENCONFIG2_DEN_RLY_CFG_RLY8_LSB = 7;
parameter DENCONFIG2_DEN_RLY_CFG_RLY8_MASK = 8'h80;
parameter DENCONFIG2_DEN_RLY_CFG_RLY8_RESET = 1'h0;


// DenConfig3
parameter DENCONFIG3_ADDR = 8'h6;
parameter DENCONFIG3_RESET = 8'h0;

// DenConfig3.DEN_DRV_CFG_RLY9
parameter DENCONFIG3_DEN_DRV_CFG_RLY9_WIDTH = 1;
parameter DENCONFIG3_DEN_DRV_CFG_RLY9_LSB = 0;
parameter DENCONFIG3_DEN_DRV_CFG_RLY9_MASK = 8'h1;
parameter DENCONFIG3_DEN_DRV_CFG_RLY9_RESET = 1'h0;

// DenConfig3.DEN_RLY_CFG_RLY9
parameter DENCONFIG3_DEN_RLY_CFG_RLY9_WIDTH = 1;
parameter DENCONFIG3_DEN_RLY_CFG_RLY9_LSB = 1;
parameter DENCONFIG3_DEN_RLY_CFG_RLY9_MASK = 8'h2;
parameter DENCONFIG3_DEN_RLY_CFG_RLY9_RESET = 1'h0;

// DenConfig3.DEN_DRV_CFG_VLV1
parameter DENCONFIG3_DEN_DRV_CFG_VLV1_WIDTH = 1;
parameter DENCONFIG3_DEN_DRV_CFG_VLV1_LSB = 2;
parameter DENCONFIG3_DEN_DRV_CFG_VLV1_MASK = 8'h4;
parameter DENCONFIG3_DEN_DRV_CFG_VLV1_RESET = 1'h0;

// DenConfig3.DEN_RLY_CFG_VLV1
parameter DENCONFIG3_DEN_RLY_CFG_VLV1_WIDTH = 1;
parameter DENCONFIG3_DEN_RLY_CFG_VLV1_LSB = 3;
parameter DENCONFIG3_DEN_RLY_CFG_VLV1_MASK = 8'h8;
parameter DENCONFIG3_DEN_RLY_CFG_VLV1_RESET = 1'h0;

// DenConfig3.DEN_DRV_CFG_VLV2
parameter DENCONFIG3_DEN_DRV_CFG_VLV2_WIDTH = 1;
parameter DENCONFIG3_DEN_DRV_CFG_VLV2_LSB = 4;
parameter DENCONFIG3_DEN_DRV_CFG_VLV2_MASK = 8'h10;
parameter DENCONFIG3_DEN_DRV_CFG_VLV2_RESET = 1'h0;

// DenConfig3.DEN_RLY_CFG_VLV2
parameter DENCONFIG3_DEN_RLY_CFG_VLV2_WIDTH = 1;
parameter DENCONFIG3_DEN_RLY_CFG_VLV2_LSB = 5;
parameter DENCONFIG3_DEN_RLY_CFG_VLV2_MASK = 8'h20;
parameter DENCONFIG3_DEN_RLY_CFG_VLV2_RESET = 1'h0;

// DenConfig3.DEN_DRV_CFG_VLV3
parameter DENCONFIG3_DEN_DRV_CFG_VLV3_WIDTH = 1;
parameter DENCONFIG3_DEN_DRV_CFG_VLV3_LSB = 6;
parameter DENCONFIG3_DEN_DRV_CFG_VLV3_MASK = 8'h40;
parameter DENCONFIG3_DEN_DRV_CFG_VLV3_RESET = 1'h0;

// DenConfig3.DEN_RLY_CFG_VLV3
parameter DENCONFIG3_DEN_RLY_CFG_VLV3_WIDTH = 1;
parameter DENCONFIG3_DEN_RLY_CFG_VLV3_LSB = 7;
parameter DENCONFIG3_DEN_RLY_CFG_VLV3_MASK = 8'h80;
parameter DENCONFIG3_DEN_RLY_CFG_VLV3_RESET = 1'h0;


// DenConfig4
parameter DENCONFIG4_ADDR = 8'h7;
parameter DENCONFIG4_RESET = 8'h0;

// DenConfig4.DEN_DRV_CFG_HTR1
parameter DENCONFIG4_DEN_DRV_CFG_HTR1_WIDTH = 1;
parameter DENCONFIG4_DEN_DRV_CFG_HTR1_LSB = 0;
parameter DENCONFIG4_DEN_DRV_CFG_HTR1_MASK = 8'h1;
parameter DENCONFIG4_DEN_DRV_CFG_HTR1_RESET = 1'h0;

// DenConfig4.DEN_RLY_CFG_HTR1
parameter DENCONFIG4_DEN_RLY_CFG_HTR1_WIDTH = 1;
parameter DENCONFIG4_DEN_RLY_CFG_HTR1_LSB = 1;
parameter DENCONFIG4_DEN_RLY_CFG_HTR1_MASK = 8'h2;
parameter DENCONFIG4_DEN_RLY_CFG_HTR1_RESET = 1'h0;

// DenConfig4.DEN_DRV_CFG_HTR2
parameter DENCONFIG4_DEN_DRV_CFG_HTR2_WIDTH = 1;
parameter DENCONFIG4_DEN_DRV_CFG_HTR2_LSB = 2;
parameter DENCONFIG4_DEN_DRV_CFG_HTR2_MASK = 8'h4;
parameter DENCONFIG4_DEN_DRV_CFG_HTR2_RESET = 1'h0;

// DenConfig4.DEN_RLY_CFG_HTR2
parameter DENCONFIG4_DEN_RLY_CFG_HTR2_WIDTH = 1;
parameter DENCONFIG4_DEN_RLY_CFG_HTR2_LSB = 3;
parameter DENCONFIG4_DEN_RLY_CFG_HTR2_MASK = 8'h8;
parameter DENCONFIG4_DEN_RLY_CFG_HTR2_RESET = 1'h0;

// DenConfig4.DEN_DRV_CFG_HB1
parameter DENCONFIG4_DEN_DRV_CFG_HB1_WIDTH = 1;
parameter DENCONFIG4_DEN_DRV_CFG_HB1_LSB = 4;
parameter DENCONFIG4_DEN_DRV_CFG_HB1_MASK = 8'h10;
parameter DENCONFIG4_DEN_DRV_CFG_HB1_RESET = 1'h0;

// DenConfig4.DEN_RLY_CFG_HB1
parameter DENCONFIG4_DEN_RLY_CFG_HB1_WIDTH = 1;
parameter DENCONFIG4_DEN_RLY_CFG_HB1_LSB = 5;
parameter DENCONFIG4_DEN_RLY_CFG_HB1_MASK = 8'h20;
parameter DENCONFIG4_DEN_RLY_CFG_HB1_RESET = 1'h0;

// DenConfig4.DEN_DRV_CFG_HB2
parameter DENCONFIG4_DEN_DRV_CFG_HB2_WIDTH = 1;
parameter DENCONFIG4_DEN_DRV_CFG_HB2_LSB = 6;
parameter DENCONFIG4_DEN_DRV_CFG_HB2_MASK = 8'h40;
parameter DENCONFIG4_DEN_DRV_CFG_HB2_RESET = 1'h0;

// DenConfig4.DEN_RLY_CFG_HB2
parameter DENCONFIG4_DEN_RLY_CFG_HB2_WIDTH = 1;
parameter DENCONFIG4_DEN_RLY_CFG_HB2_LSB = 7;
parameter DENCONFIG4_DEN_RLY_CFG_HB2_MASK = 8'h80;
parameter DENCONFIG4_DEN_RLY_CFG_HB2_RESET = 1'h0;


// OEConfig0
parameter OECONFIG0_ADDR = 8'h8;
parameter OECONFIG0_RESET = 8'h0;

// OEConfig0.IGN_OE
parameter OECONFIG0_IGN_OE_WIDTH = 4;
parameter OECONFIG0_IGN_OE_LSB = 0;
parameter OECONFIG0_IGN_OE_MASK = 8'hf;
parameter OECONFIG0_IGN_OE_RESET = 4'h0;

// OEConfig0.INJ_OE
parameter OECONFIG0_INJ_OE_WIDTH = 4;
parameter OECONFIG0_INJ_OE_LSB = 4;
parameter OECONFIG0_INJ_OE_MASK = 8'hf0;
parameter OECONFIG0_INJ_OE_RESET = 4'h0;


// OEConfig1
parameter OECONFIG1_ADDR = 8'h9;
parameter OECONFIG1_RESET = 8'h0;

// OEConfig1.RLY_OE
parameter OECONFIG1_RLY_OE_WIDTH = 8;
parameter OECONFIG1_RLY_OE_LSB = 0;
parameter OECONFIG1_RLY_OE_MASK = 8'hff;
parameter OECONFIG1_RLY_OE_RESET = 8'h0;


// OEConfig2
parameter OECONFIG2_ADDR = 8'ha;
parameter OECONFIG2_RESET = 8'h0;

// OEConfig2.RLY_OE
parameter OECONFIG2_RLY_OE_WIDTH = 1;
parameter OECONFIG2_RLY_OE_LSB = 0;
parameter OECONFIG2_RLY_OE_MASK = 8'h1;
parameter OECONFIG2_RLY_OE_RESET = 1'h0;

// OEConfig2.HTR_OE
parameter OECONFIG2_HTR_OE_WIDTH = 2;
parameter OECONFIG2_HTR_OE_LSB = 1;
parameter OECONFIG2_HTR_OE_MASK = 8'h6;
parameter OECONFIG2_HTR_OE_RESET = 2'h0;

// OEConfig2.VLV_OE
parameter OECONFIG2_VLV_OE_WIDTH = 3;
parameter OECONFIG2_VLV_OE_LSB = 3;
parameter OECONFIG2_VLV_OE_MASK = 8'h38;
parameter OECONFIG2_VLV_OE_RESET = 3'h0;


// OEConfig3
parameter OECONFIG3_ADDR = 8'hb;
parameter OECONFIG3_RESET = 8'h0;

// OEConfig3.HS_OE
parameter OECONFIG3_HS_OE_WIDTH = 2;
parameter OECONFIG3_HS_OE_LSB = 0;
parameter OECONFIG3_HS_OE_MASK = 8'h3;
parameter OECONFIG3_HS_OE_RESET = 2'h0;

// OEConfig3.LS_OE
parameter OECONFIG3_LS_OE_WIDTH = 2;
parameter OECONFIG3_LS_OE_LSB = 2;
parameter OECONFIG3_LS_OE_MASK = 8'hc;
parameter OECONFIG3_LS_OE_RESET = 2'h0;


// DDConfig0
parameter DDCONFIG0_ADDR = 8'hc;
parameter DDCONFIG0_RESET = 8'h0;

// DDConfig0.IGN_DD
parameter DDCONFIG0_IGN_DD_WIDTH = 4;
parameter DDCONFIG0_IGN_DD_LSB = 0;
parameter DDCONFIG0_IGN_DD_MASK = 8'hf;
parameter DDCONFIG0_IGN_DD_RESET = 4'h0;

// DDConfig0.INJ_DD
parameter DDCONFIG0_INJ_DD_WIDTH = 4;
parameter DDCONFIG0_INJ_DD_LSB = 4;
parameter DDCONFIG0_INJ_DD_MASK = 8'hf0;
parameter DDCONFIG0_INJ_DD_RESET = 4'h0;


// DDConfig1
parameter DDCONFIG1_ADDR = 8'hd;
parameter DDCONFIG1_RESET = 8'h0;

// DDConfig1.RLY_DD
parameter DDCONFIG1_RLY_DD_WIDTH = 8;
parameter DDCONFIG1_RLY_DD_LSB = 0;
parameter DDCONFIG1_RLY_DD_MASK = 8'hff;
parameter DDCONFIG1_RLY_DD_RESET = 8'h0;


// DDConfig2
parameter DDCONFIG2_ADDR = 8'he;
parameter DDCONFIG2_RESET = 8'h0;

// DDConfig2.RLY_DD
parameter DDCONFIG2_RLY_DD_WIDTH = 1;
parameter DDCONFIG2_RLY_DD_LSB = 0;
parameter DDCONFIG2_RLY_DD_MASK = 8'h1;
parameter DDCONFIG2_RLY_DD_RESET = 1'h0;

// DDConfig2.HTR_DD
parameter DDCONFIG2_HTR_DD_WIDTH = 2;
parameter DDCONFIG2_HTR_DD_LSB = 1;
parameter DDCONFIG2_HTR_DD_MASK = 8'h6;
parameter DDCONFIG2_HTR_DD_RESET = 2'h0;

// DDConfig2.VLV_DD
parameter DDCONFIG2_VLV_DD_WIDTH = 3;
parameter DDCONFIG2_VLV_DD_LSB = 3;
parameter DDCONFIG2_VLV_DD_MASK = 8'h38;
parameter DDCONFIG2_VLV_DD_RESET = 3'h0;

// DDConfig2.HB_DD
parameter DDCONFIG2_HB_DD_WIDTH = 2;
parameter DDCONFIG2_HB_DD_LSB = 6;
parameter DDCONFIG2_HB_DD_MASK = 8'hc0;
parameter DDCONFIG2_HB_DD_RESET = 2'h0;


// Cont0
parameter CONT0_ADDR = 8'hf;
parameter CONT0_RESET = 8'h0;

// Cont0.IGN_ON
parameter CONT0_IGN_ON_WIDTH = 4;
parameter CONT0_IGN_ON_LSB = 0;
parameter CONT0_IGN_ON_MASK = 8'hf;
parameter CONT0_IGN_ON_RESET = 4'h0;

// Cont0.INJ_ON
parameter CONT0_INJ_ON_WIDTH = 4;
parameter CONT0_INJ_ON_LSB = 4;
parameter CONT0_INJ_ON_MASK = 8'hf0;
parameter CONT0_INJ_ON_RESET = 4'h0;


// Cont1
parameter CONT1_ADDR = 8'h10;
parameter CONT1_RESET = 8'h0;

// Cont1.RLY_ON
parameter CONT1_RLY_ON_WIDTH = 8;
parameter CONT1_RLY_ON_LSB = 0;
parameter CONT1_RLY_ON_MASK = 8'hff;
parameter CONT1_RLY_ON_RESET = 8'h0;


// Cont2
parameter CONT2_ADDR = 8'h11;
parameter CONT2_RESET = 8'h0;

// Cont2.RLY_ON
parameter CONT2_RLY_ON_WIDTH = 1;
parameter CONT2_RLY_ON_LSB = 0;
parameter CONT2_RLY_ON_MASK = 8'h1;
parameter CONT2_RLY_ON_RESET = 1'h0;

// Cont2.HTR_ON
parameter CONT2_HTR_ON_WIDTH = 2;
parameter CONT2_HTR_ON_LSB = 1;
parameter CONT2_HTR_ON_MASK = 8'h6;
parameter CONT2_HTR_ON_RESET = 2'h0;

// Cont2.VLV_ON
parameter CONT2_VLV_ON_WIDTH = 3;
parameter CONT2_VLV_ON_LSB = 3;
parameter CONT2_VLV_ON_MASK = 8'h38;
parameter CONT2_VLV_ON_RESET = 3'h0;

// Cont2.HB_ON
parameter CONT2_HB_ON_WIDTH = 2;
parameter CONT2_HB_ON_LSB = 6;
parameter CONT2_HB_ON_MASK = 8'hc0;
parameter CONT2_HB_ON_RESET = 2'h0;


// BRIConfig0
parameter BRICONFIG0_ADDR = 8'h12;
parameter BRICONFIG0_RESET = 8'h0;

// BRIConfig0.FW_MODE
parameter BRICONFIG0_FW_MODE_WIDTH = 2;
parameter BRICONFIG0_FW_MODE_LSB = 0;
parameter BRICONFIG0_FW_MODE_MASK = 8'h3;
parameter BRICONFIG0_FW_MODE_RESET = 2'h0;

// BRIConfig0.HS_LS_MODE
parameter BRICONFIG0_HS_LS_MODE_WIDTH = 2;
parameter BRICONFIG0_HS_LS_MODE_LSB = 2;
parameter BRICONFIG0_HS_LS_MODE_MASK = 8'hc;
parameter BRICONFIG0_HS_LS_MODE_RESET = 2'h0;


// IgnDiagConfig
parameter IGNDIAGCONFIG_ADDR = 8'h13;
parameter IGNDIAGCONFIG_RESET = 8'h5;

// IgnDiagConfig.EN_DIAG_OL_IGN
parameter IGNDIAGCONFIG_EN_DIAG_OL_IGN_WIDTH = 1;
parameter IGNDIAGCONFIG_EN_DIAG_OL_IGN_LSB = 0;
parameter IGNDIAGCONFIG_EN_DIAG_OL_IGN_MASK = 8'h1;
parameter IGNDIAGCONFIG_EN_DIAG_OL_IGN_RESET = 1'h1;

// IgnDiagConfig.SEL_OL_TH_IGN
parameter IGNDIAGCONFIG_SEL_OL_TH_IGN_WIDTH = 2;
parameter IGNDIAGCONFIG_SEL_OL_TH_IGN_LSB = 1;
parameter IGNDIAGCONFIG_SEL_OL_TH_IGN_MASK = 8'h6;
parameter IGNDIAGCONFIG_SEL_OL_TH_IGN_RESET = 2'h2;


// OutDiagConfig0
parameter OUTDIAGCONFIG0_ADDR = 8'h14;
parameter OUTDIAGCONFIG0_RESET = 8'hff;

// OutDiagConfig0.DIAG_INJ1
parameter OUTDIAGCONFIG0_DIAG_INJ1_WIDTH = 2;
parameter OUTDIAGCONFIG0_DIAG_INJ1_LSB = 0;
parameter OUTDIAGCONFIG0_DIAG_INJ1_MASK = 8'h3;
parameter OUTDIAGCONFIG0_DIAG_INJ1_RESET = 2'h3;

// OutDiagConfig0.DIAG_INJ2
parameter OUTDIAGCONFIG0_DIAG_INJ2_WIDTH = 2;
parameter OUTDIAGCONFIG0_DIAG_INJ2_LSB = 2;
parameter OUTDIAGCONFIG0_DIAG_INJ2_MASK = 8'hc;
parameter OUTDIAGCONFIG0_DIAG_INJ2_RESET = 2'h3;

// OutDiagConfig0.DIAG_INJ3
parameter OUTDIAGCONFIG0_DIAG_INJ3_WIDTH = 2;
parameter OUTDIAGCONFIG0_DIAG_INJ3_LSB = 4;
parameter OUTDIAGCONFIG0_DIAG_INJ3_MASK = 8'h30;
parameter OUTDIAGCONFIG0_DIAG_INJ3_RESET = 2'h3;

// OutDiagConfig0.DIAG_INJ4
parameter OUTDIAGCONFIG0_DIAG_INJ4_WIDTH = 2;
parameter OUTDIAGCONFIG0_DIAG_INJ4_LSB = 6;
parameter OUTDIAGCONFIG0_DIAG_INJ4_MASK = 8'hc0;
parameter OUTDIAGCONFIG0_DIAG_INJ4_RESET = 2'h3;


// OutDiagConfig1
parameter OUTDIAGCONFIG1_ADDR = 8'h15;
parameter OUTDIAGCONFIG1_RESET = 8'hff;

// OutDiagConfig1.DIAG_RLY1
parameter OUTDIAGCONFIG1_DIAG_RLY1_WIDTH = 2;
parameter OUTDIAGCONFIG1_DIAG_RLY1_LSB = 0;
parameter OUTDIAGCONFIG1_DIAG_RLY1_MASK = 8'h3;
parameter OUTDIAGCONFIG1_DIAG_RLY1_RESET = 2'h3;

// OutDiagConfig1.DIAG_RLY2
parameter OUTDIAGCONFIG1_DIAG_RLY2_WIDTH = 2;
parameter OUTDIAGCONFIG1_DIAG_RLY2_LSB = 2;
parameter OUTDIAGCONFIG1_DIAG_RLY2_MASK = 8'hc;
parameter OUTDIAGCONFIG1_DIAG_RLY2_RESET = 2'h3;

// OutDiagConfig1.DIAG_RLY3
parameter OUTDIAGCONFIG1_DIAG_RLY3_WIDTH = 2;
parameter OUTDIAGCONFIG1_DIAG_RLY3_LSB = 4;
parameter OUTDIAGCONFIG1_DIAG_RLY3_MASK = 8'h30;
parameter OUTDIAGCONFIG1_DIAG_RLY3_RESET = 2'h3;

// OutDiagConfig1.DIAG_RLY4
parameter OUTDIAGCONFIG1_DIAG_RLY4_WIDTH = 2;
parameter OUTDIAGCONFIG1_DIAG_RLY4_LSB = 6;
parameter OUTDIAGCONFIG1_DIAG_RLY4_MASK = 8'hc0;
parameter OUTDIAGCONFIG1_DIAG_RLY4_RESET = 2'h3;


// OutDiagConfig2
parameter OUTDIAGCONFIG2_ADDR = 8'h16;
parameter OUTDIAGCONFIG2_RESET = 8'hff;

// OutDiagConfig2.DIAG_RLY5
parameter OUTDIAGCONFIG2_DIAG_RLY5_WIDTH = 2;
parameter OUTDIAGCONFIG2_DIAG_RLY5_LSB = 0;
parameter OUTDIAGCONFIG2_DIAG_RLY5_MASK = 8'h3;
parameter OUTDIAGCONFIG2_DIAG_RLY5_RESET = 2'h3;

// OutDiagConfig2.DIAG_RLY6
parameter OUTDIAGCONFIG2_DIAG_RLY6_WIDTH = 2;
parameter OUTDIAGCONFIG2_DIAG_RLY6_LSB = 2;
parameter OUTDIAGCONFIG2_DIAG_RLY6_MASK = 8'hc;
parameter OUTDIAGCONFIG2_DIAG_RLY6_RESET = 2'h3;

// OutDiagConfig2.DIAG_RLY7
parameter OUTDIAGCONFIG2_DIAG_RLY7_WIDTH = 2;
parameter OUTDIAGCONFIG2_DIAG_RLY7_LSB = 4;
parameter OUTDIAGCONFIG2_DIAG_RLY7_MASK = 8'h30;
parameter OUTDIAGCONFIG2_DIAG_RLY7_RESET = 2'h3;

// OutDiagConfig2.DIAG_RLY8
parameter OUTDIAGCONFIG2_DIAG_RLY8_WIDTH = 2;
parameter OUTDIAGCONFIG2_DIAG_RLY8_LSB = 6;
parameter OUTDIAGCONFIG2_DIAG_RLY8_MASK = 8'hc0;
parameter OUTDIAGCONFIG2_DIAG_RLY8_RESET = 2'h3;


// OutDiagConfig3
parameter OUTDIAGCONFIG3_ADDR = 8'h17;
parameter OUTDIAGCONFIG3_RESET = 8'hff;

// OutDiagConfig3.DIAG_RLY9
parameter OUTDIAGCONFIG3_DIAG_RLY9_WIDTH = 2;
parameter OUTDIAGCONFIG3_DIAG_RLY9_LSB = 0;
parameter OUTDIAGCONFIG3_DIAG_RLY9_MASK = 8'h3;
parameter OUTDIAGCONFIG3_DIAG_RLY9_RESET = 2'h3;

// OutDiagConfig3.DIAG_VLV1
parameter OUTDIAGCONFIG3_DIAG_VLV1_WIDTH = 2;
parameter OUTDIAGCONFIG3_DIAG_VLV1_LSB = 2;
parameter OUTDIAGCONFIG3_DIAG_VLV1_MASK = 8'hc;
parameter OUTDIAGCONFIG3_DIAG_VLV1_RESET = 2'h3;

// OutDiagConfig3.DIAG_VLV2
parameter OUTDIAGCONFIG3_DIAG_VLV2_WIDTH = 2;
parameter OUTDIAGCONFIG3_DIAG_VLV2_LSB = 4;
parameter OUTDIAGCONFIG3_DIAG_VLV2_MASK = 8'h30;
parameter OUTDIAGCONFIG3_DIAG_VLV2_RESET = 2'h3;

// OutDiagConfig3.DIAG_VLV3
parameter OUTDIAGCONFIG3_DIAG_VLV3_WIDTH = 2;
parameter OUTDIAGCONFIG3_DIAG_VLV3_LSB = 6;
parameter OUTDIAGCONFIG3_DIAG_VLV3_MASK = 8'hc0;
parameter OUTDIAGCONFIG3_DIAG_VLV3_RESET = 2'h3;


// OutDiagConfig4
parameter OUTDIAGCONFIG4_ADDR = 8'h18;
parameter OUTDIAGCONFIG4_RESET = 8'hff;

// OutDiagConfig4.DIAG_HTR1
parameter OUTDIAGCONFIG4_DIAG_HTR1_WIDTH = 2;
parameter OUTDIAGCONFIG4_DIAG_HTR1_LSB = 0;
parameter OUTDIAGCONFIG4_DIAG_HTR1_MASK = 8'h3;
parameter OUTDIAGCONFIG4_DIAG_HTR1_RESET = 2'h3;

// OutDiagConfig4.DIAG_HTR2
parameter OUTDIAGCONFIG4_DIAG_HTR2_WIDTH = 2;
parameter OUTDIAGCONFIG4_DIAG_HTR2_LSB = 2;
parameter OUTDIAGCONFIG4_DIAG_HTR2_MASK = 8'hc;
parameter OUTDIAGCONFIG4_DIAG_HTR2_RESET = 2'h3;

// OutDiagConfig4.DIAG_HB1
parameter OUTDIAGCONFIG4_DIAG_HB1_WIDTH = 2;
parameter OUTDIAGCONFIG4_DIAG_HB1_LSB = 4;
parameter OUTDIAGCONFIG4_DIAG_HB1_MASK = 8'h30;
parameter OUTDIAGCONFIG4_DIAG_HB1_RESET = 2'h3;

// OutDiagConfig4.DIAG_HB2
parameter OUTDIAGCONFIG4_DIAG_HB2_WIDTH = 2;
parameter OUTDIAGCONFIG4_DIAG_HB2_LSB = 6;
parameter OUTDIAGCONFIG4_DIAG_HB2_MASK = 8'hc0;
parameter OUTDIAGCONFIG4_DIAG_HB2_RESET = 2'h3;


// CurrLimConfig0
parameter CURRLIMCONFIG0_ADDR = 8'h19;
parameter CURRLIMCONFIG0_RESET = 8'h0;

// CurrLimConfig0.CURR_LIM_INJ
parameter CURRLIMCONFIG0_CURR_LIM_INJ_WIDTH = 4;
parameter CURRLIMCONFIG0_CURR_LIM_INJ_LSB = 0;
parameter CURRLIMCONFIG0_CURR_LIM_INJ_MASK = 8'hf;
parameter CURRLIMCONFIG0_CURR_LIM_INJ_RESET = 4'h0;


// CurrLimConfig1
parameter CURRLIMCONFIG1_ADDR = 8'h1a;
parameter CURRLIMCONFIG1_RESET = 8'h0;

// CurrLimConfig1.CURR_LIM_RLY
parameter CURRLIMCONFIG1_CURR_LIM_RLY_WIDTH = 8;
parameter CURRLIMCONFIG1_CURR_LIM_RLY_LSB = 0;
parameter CURRLIMCONFIG1_CURR_LIM_RLY_MASK = 8'hff;
parameter CURRLIMCONFIG1_CURR_LIM_RLY_RESET = 8'h0;


// CurrLimConfig2
parameter CURRLIMCONFIG2_ADDR = 8'h1b;
parameter CURRLIMCONFIG2_RESET = 8'h0;

// CurrLimConfig2.CURR_LIM_RLY
parameter CURRLIMCONFIG2_CURR_LIM_RLY_WIDTH = 1;
parameter CURRLIMCONFIG2_CURR_LIM_RLY_LSB = 0;
parameter CURRLIMCONFIG2_CURR_LIM_RLY_MASK = 8'h1;
parameter CURRLIMCONFIG2_CURR_LIM_RLY_RESET = 1'h0;

// CurrLimConfig2.CURR_LIM_VLV
parameter CURRLIMCONFIG2_CURR_LIM_VLV_WIDTH = 3;
parameter CURRLIMCONFIG2_CURR_LIM_VLV_LSB = 1;
parameter CURRLIMCONFIG2_CURR_LIM_VLV_MASK = 8'he;
parameter CURRLIMCONFIG2_CURR_LIM_VLV_RESET = 3'h0;

// CurrLimConfig2.CURR_LIM_HTR
parameter CURRLIMCONFIG2_CURR_LIM_HTR_WIDTH = 2;
parameter CURRLIMCONFIG2_CURR_LIM_HTR_LSB = 4;
parameter CURRLIMCONFIG2_CURR_LIM_HTR_MASK = 8'h30;
parameter CURRLIMCONFIG2_CURR_LIM_HTR_RESET = 2'h0;

// CurrLimConfig2.CURR_LIM_HB
parameter CURRLIMCONFIG2_CURR_LIM_HB_WIDTH = 2;
parameter CURRLIMCONFIG2_CURR_LIM_HB_LSB = 6;
parameter CURRLIMCONFIG2_CURR_LIM_HB_MASK = 8'hc0;
parameter CURRLIMCONFIG2_CURR_LIM_HB_RESET = 2'h0;


// DlyOffConfig
parameter DLYOFFCONFIG_ADDR = 8'h1c;
parameter DLYOFFCONFIG_RESET = 8'h0;

// DlyOffConfig.DEL_OFF_RLY
parameter DLYOFFCONFIG_DEL_OFF_RLY_WIDTH = 3;
parameter DLYOFFCONFIG_DEL_OFF_RLY_LSB = 0;
parameter DLYOFFCONFIG_DEL_OFF_RLY_MASK = 8'h7;
parameter DLYOFFCONFIG_DEL_OFF_RLY_RESET = 3'h0;

// DlyOffConfig.DEL_OFF_HB
parameter DLYOFFCONFIG_DEL_OFF_HB_WIDTH = 2;
parameter DLYOFFCONFIG_DEL_OFF_HB_LSB = 3;
parameter DLYOFFCONFIG_DEL_OFF_HB_MASK = 8'h18;
parameter DLYOFFCONFIG_DEL_OFF_HB_RESET = 2'h0;


// DinConfig0
parameter DINCONFIG0_ADDR = 8'h1d;
parameter DINCONFIG0_RESET = 8'h21;

// DinConfig0.INJ_IN1
parameter DINCONFIG0_INJ_IN1_WIDTH = 4;
parameter DINCONFIG0_INJ_IN1_LSB = 0;
parameter DINCONFIG0_INJ_IN1_MASK = 8'hf;
parameter DINCONFIG0_INJ_IN1_RESET = 4'h1;

// DinConfig0.INJ_IN2
parameter DINCONFIG0_INJ_IN2_WIDTH = 4;
parameter DINCONFIG0_INJ_IN2_LSB = 4;
parameter DINCONFIG0_INJ_IN2_MASK = 8'hf0;
parameter DINCONFIG0_INJ_IN2_RESET = 4'h2;


// DinConfig1
parameter DINCONFIG1_ADDR = 8'h1e;
parameter DINCONFIG1_RESET = 8'h43;

// DinConfig1.INJ_IN3
parameter DINCONFIG1_INJ_IN3_WIDTH = 4;
parameter DINCONFIG1_INJ_IN3_LSB = 0;
parameter DINCONFIG1_INJ_IN3_MASK = 8'hf;
parameter DINCONFIG1_INJ_IN3_RESET = 4'h3;

// DinConfig1.INJ_IN4
parameter DINCONFIG1_INJ_IN4_WIDTH = 4;
parameter DINCONFIG1_INJ_IN4_LSB = 4;
parameter DINCONFIG1_INJ_IN4_MASK = 8'hf0;
parameter DINCONFIG1_INJ_IN4_RESET = 4'h4;


// DinConfig2
parameter DINCONFIG2_ADDR = 8'h1f;
parameter DINCONFIG2_RESET = 8'hba;

// DinConfig2.IGN_IN1
parameter DINCONFIG2_IGN_IN1_WIDTH = 4;
parameter DINCONFIG2_IGN_IN1_LSB = 0;
parameter DINCONFIG2_IGN_IN1_MASK = 8'hf;
parameter DINCONFIG2_IGN_IN1_RESET = 4'ha;

// DinConfig2.IGN_IN2
parameter DINCONFIG2_IGN_IN2_WIDTH = 4;
parameter DINCONFIG2_IGN_IN2_LSB = 4;
parameter DINCONFIG2_IGN_IN2_MASK = 8'hf0;
parameter DINCONFIG2_IGN_IN2_RESET = 4'hb;


// DinConfig3
parameter DINCONFIG3_ADDR = 8'h20;
parameter DINCONFIG3_RESET = 8'hdc;

// DinConfig3.IGN_IN3
parameter DINCONFIG3_IGN_IN3_WIDTH = 4;
parameter DINCONFIG3_IGN_IN3_LSB = 0;
parameter DINCONFIG3_IGN_IN3_MASK = 8'hf;
parameter DINCONFIG3_IGN_IN3_RESET = 4'hc;

// DinConfig3.IGN_IN4
parameter DINCONFIG3_IGN_IN4_WIDTH = 4;
parameter DINCONFIG3_IGN_IN4_LSB = 4;
parameter DINCONFIG3_IGN_IN4_MASK = 8'hf0;
parameter DINCONFIG3_IGN_IN4_RESET = 4'hd;


// DinConfig4
parameter DINCONFIG4_ADDR = 8'h21;
parameter DINCONFIG4_RESET = 8'h0;

// DinConfig4.HTR_IN1
parameter DINCONFIG4_HTR_IN1_WIDTH = 4;
parameter DINCONFIG4_HTR_IN1_LSB = 0;
parameter DINCONFIG4_HTR_IN1_MASK = 8'hf;
parameter DINCONFIG4_HTR_IN1_RESET = 4'h0;

// DinConfig4.HTR_IN2
parameter DINCONFIG4_HTR_IN2_WIDTH = 4;
parameter DINCONFIG4_HTR_IN2_LSB = 4;
parameter DINCONFIG4_HTR_IN2_MASK = 8'hf0;
parameter DINCONFIG4_HTR_IN2_RESET = 4'h0;


// DinConfig5
parameter DINCONFIG5_ADDR = 8'h22;
parameter DINCONFIG5_RESET = 8'h0;

// DinConfig5.HB_IN1
parameter DINCONFIG5_HB_IN1_WIDTH = 4;
parameter DINCONFIG5_HB_IN1_LSB = 0;
parameter DINCONFIG5_HB_IN1_MASK = 8'hf;
parameter DINCONFIG5_HB_IN1_RESET = 4'h0;

// DinConfig5.HB_IN2
parameter DINCONFIG5_HB_IN2_WIDTH = 4;
parameter DINCONFIG5_HB_IN2_LSB = 4;
parameter DINCONFIG5_HB_IN2_MASK = 8'hf0;
parameter DINCONFIG5_HB_IN2_RESET = 4'h0;


// DinConfig6
parameter DINCONFIG6_ADDR = 8'h23;
parameter DINCONFIG6_RESET = 8'h0;

// DinConfig6.RLY_IN1
parameter DINCONFIG6_RLY_IN1_WIDTH = 4;
parameter DINCONFIG6_RLY_IN1_LSB = 0;
parameter DINCONFIG6_RLY_IN1_MASK = 8'hf;
parameter DINCONFIG6_RLY_IN1_RESET = 4'h0;

// DinConfig6.RLY_IN2
parameter DINCONFIG6_RLY_IN2_WIDTH = 4;
parameter DINCONFIG6_RLY_IN2_LSB = 4;
parameter DINCONFIG6_RLY_IN2_MASK = 8'hf0;
parameter DINCONFIG6_RLY_IN2_RESET = 4'h0;


// DinConfig7
parameter DINCONFIG7_ADDR = 8'h24;
parameter DINCONFIG7_RESET = 8'h0;

// DinConfig7.RLY_IN3
parameter DINCONFIG7_RLY_IN3_WIDTH = 4;
parameter DINCONFIG7_RLY_IN3_LSB = 0;
parameter DINCONFIG7_RLY_IN3_MASK = 8'hf;
parameter DINCONFIG7_RLY_IN3_RESET = 4'h0;

// DinConfig7.RLY_IN4
parameter DINCONFIG7_RLY_IN4_WIDTH = 4;
parameter DINCONFIG7_RLY_IN4_LSB = 4;
parameter DINCONFIG7_RLY_IN4_MASK = 8'hf0;
parameter DINCONFIG7_RLY_IN4_RESET = 4'h0;


// DinConfig8
parameter DINCONFIG8_ADDR = 8'h25;
parameter DINCONFIG8_RESET = 8'h0;

// DinConfig8.RLY_IN5
parameter DINCONFIG8_RLY_IN5_WIDTH = 4;
parameter DINCONFIG8_RLY_IN5_LSB = 0;
parameter DINCONFIG8_RLY_IN5_MASK = 8'hf;
parameter DINCONFIG8_RLY_IN5_RESET = 4'h0;

// DinConfig8.RLY_IN6
parameter DINCONFIG8_RLY_IN6_WIDTH = 4;
parameter DINCONFIG8_RLY_IN6_LSB = 4;
parameter DINCONFIG8_RLY_IN6_MASK = 8'hf0;
parameter DINCONFIG8_RLY_IN6_RESET = 4'h0;


// DinConfig9
parameter DINCONFIG9_ADDR = 8'h26;
parameter DINCONFIG9_RESET = 8'h80;

// DinConfig9.RLY_IN7
parameter DINCONFIG9_RLY_IN7_WIDTH = 4;
parameter DINCONFIG9_RLY_IN7_LSB = 0;
parameter DINCONFIG9_RLY_IN7_MASK = 8'hf;
parameter DINCONFIG9_RLY_IN7_RESET = 4'h0;

// DinConfig9.RLY_IN8
parameter DINCONFIG9_RLY_IN8_WIDTH = 4;
parameter DINCONFIG9_RLY_IN8_LSB = 4;
parameter DINCONFIG9_RLY_IN8_MASK = 8'hf0;
parameter DINCONFIG9_RLY_IN8_RESET = 4'h8;


// DinConfig10
parameter DINCONFIG10_ADDR = 8'h27;
parameter DINCONFIG10_RESET = 8'h59;

// DinConfig10.RLY_IN9
parameter DINCONFIG10_RLY_IN9_WIDTH = 4;
parameter DINCONFIG10_RLY_IN9_LSB = 0;
parameter DINCONFIG10_RLY_IN9_MASK = 8'hf;
parameter DINCONFIG10_RLY_IN9_RESET = 4'h9;

// DinConfig10.VLV_IN1
parameter DINCONFIG10_VLV_IN1_WIDTH = 4;
parameter DINCONFIG10_VLV_IN1_LSB = 4;
parameter DINCONFIG10_VLV_IN1_MASK = 8'hf0;
parameter DINCONFIG10_VLV_IN1_RESET = 4'h5;


// DinConfig11
parameter DINCONFIG11_ADDR = 8'h28;
parameter DINCONFIG11_RESET = 8'h76;

// DinConfig11.VLV_IN2
parameter DINCONFIG11_VLV_IN2_WIDTH = 4;
parameter DINCONFIG11_VLV_IN2_LSB = 0;
parameter DINCONFIG11_VLV_IN2_MASK = 8'hf;
parameter DINCONFIG11_VLV_IN2_RESET = 4'h6;

// DinConfig11.VLV_IN3
parameter DINCONFIG11_VLV_IN3_WIDTH = 4;
parameter DINCONFIG11_VLV_IN3_LSB = 4;
parameter DINCONFIG11_VLV_IN3_MASK = 8'hf0;
parameter DINCONFIG11_VLV_IN3_RESET = 4'h7;


// WDConfig0
parameter WDCONFIG0_ADDR = 8'h29;
parameter WDCONFIG0_RESET = 8'h20;

// WDConfig0.WD_DURATION
parameter WDCONFIG0_WD_DURATION_WIDTH = 4;
parameter WDCONFIG0_WD_DURATION_LSB = 0;
parameter WDCONFIG0_WD_DURATION_MASK = 8'hf;
parameter WDCONFIG0_WD_DURATION_RESET = 4'h0;

// WDConfig0.VRS_WD_DURATION
parameter WDCONFIG0_VRS_WD_DURATION_WIDTH = 2;
parameter WDCONFIG0_VRS_WD_DURATION_LSB = 4;
parameter WDCONFIG0_VRS_WD_DURATION_MASK = 8'h30;
parameter WDCONFIG0_VRS_WD_DURATION_RESET = 2'h2;

// WDConfig0.VRS_WD_EN
parameter WDCONFIG0_VRS_WD_EN_WIDTH = 1;
parameter WDCONFIG0_VRS_WD_EN_LSB = 6;
parameter WDCONFIG0_VRS_WD_EN_MASK = 8'h40;
parameter WDCONFIG0_VRS_WD_EN_RESET = 1'h0;


// WDConfig1
parameter WDCONFIG1_ADDR = 8'h2a;
parameter WDCONFIG1_RESET = 8'h0;

// WDConfig1.SPI_ERR_CNT_CFG
parameter WDCONFIG1_SPI_ERR_CNT_CFG_WIDTH = 2;
parameter WDCONFIG1_SPI_ERR_CNT_CFG_LSB = 0;
parameter WDCONFIG1_SPI_ERR_CNT_CFG_MASK = 8'h3;
parameter WDCONFIG1_SPI_ERR_CNT_CFG_RESET = 2'h0;

// WDConfig1.SPI_RFH_CNT_CFG
parameter WDCONFIG1_SPI_RFH_CNT_CFG_WIDTH = 2;
parameter WDCONFIG1_SPI_RFH_CNT_CFG_LSB = 2;
parameter WDCONFIG1_SPI_RFH_CNT_CFG_MASK = 8'hc;
parameter WDCONFIG1_SPI_RFH_CNT_CFG_RESET = 2'h0;

// WDConfig1.SPI_RST_ERR_FS
parameter WDCONFIG1_SPI_RST_ERR_FS_WIDTH = 1;
parameter WDCONFIG1_SPI_RST_ERR_FS_LSB = 4;
parameter WDCONFIG1_SPI_RST_ERR_FS_MASK = 8'h10;
parameter WDCONFIG1_SPI_RST_ERR_FS_RESET = 1'h0;


// VrsConfig0
parameter VRSCONFIG0_ADDR = 8'h2b;
parameter VRSCONFIG0_RESET = 8'h2;

// VrsConfig0.VRS_MODE_CFG
parameter VRSCONFIG0_VRS_MODE_CFG_WIDTH = 2;
parameter VRSCONFIG0_VRS_MODE_CFG_LSB = 0;
parameter VRSCONFIG0_VRS_MODE_CFG_MASK = 8'h3;
parameter VRSCONFIG0_VRS_MODE_CFG_RESET = 2'h2;

// VrsConfig0.VRS_REF
parameter VRSCONFIG0_VRS_REF_WIDTH = 2;
parameter VRSCONFIG0_VRS_REF_LSB = 2;
parameter VRSCONFIG0_VRS_REF_MASK = 8'hc;
parameter VRSCONFIG0_VRS_REF_RESET = 2'h0;

// VrsConfig0.VRS_TEST_CFG
parameter VRSCONFIG0_VRS_TEST_CFG_WIDTH = 2;
parameter VRSCONFIG0_VRS_TEST_CFG_LSB = 4;
parameter VRSCONFIG0_VRS_TEST_CFG_MASK = 8'h30;
parameter VRSCONFIG0_VRS_TEST_CFG_RESET = 2'h0;

// VrsConfig0.VRSO_SPI_CTRL_MODE
parameter VRSCONFIG0_VRSO_SPI_CTRL_MODE_WIDTH = 1;
parameter VRSCONFIG0_VRSO_SPI_CTRL_MODE_LSB = 6;
parameter VRSCONFIG0_VRSO_SPI_CTRL_MODE_MASK = 8'h40;
parameter VRSCONFIG0_VRSO_SPI_CTRL_MODE_RESET = 1'h0;

// VrsConfig0.VRSO_SPI_CTRL
parameter VRSCONFIG0_VRSO_SPI_CTRL_WIDTH = 1;
parameter VRSCONFIG0_VRSO_SPI_CTRL_LSB = 7;
parameter VRSCONFIG0_VRSO_SPI_CTRL_MASK = 8'h80;
parameter VRSCONFIG0_VRSO_SPI_CTRL_RESET = 1'h0;


// VrsConfig1
parameter VRSCONFIG1_ADDR = 8'h2c;
parameter VRSCONFIG1_RESET = 8'h78;

// VrsConfig1.VRSF
parameter VRSCONFIG1_VRSF_WIDTH = 3;
parameter VRSCONFIG1_VRSF_LSB = 0;
parameter VRSCONFIG1_VRSF_MASK = 8'h7;
parameter VRSCONFIG1_VRSF_RESET = 3'h0;

// VrsConfig1.VRSM
parameter VRSCONFIG1_VRSM_WIDTH = 1;
parameter VRSCONFIG1_VRSM_LSB = 3;
parameter VRSCONFIG1_VRSM_MASK = 8'h8;
parameter VRSCONFIG1_VRSM_RESET = 1'h1;

// VrsConfig1.VRSRF
parameter VRSCONFIG1_VRSRF_WIDTH = 1;
parameter VRSCONFIG1_VRSRF_LSB = 4;
parameter VRSCONFIG1_VRSRF_MASK = 8'h10;
parameter VRSCONFIG1_VRSRF_RESET = 1'h1;

// VrsConfig1.VRSFF
parameter VRSCONFIG1_VRSFF_WIDTH = 1;
parameter VRSCONFIG1_VRSFF_LSB = 5;
parameter VRSCONFIG1_VRSFF_MASK = 8'h20;
parameter VRSCONFIG1_VRSFF_RESET = 1'h1;

// VrsConfig1.VRSEFF
parameter VRSCONFIG1_VRSEFF_WIDTH = 1;
parameter VRSCONFIG1_VRSEFF_LSB = 6;
parameter VRSCONFIG1_VRSEFF_MASK = 8'h40;
parameter VRSCONFIG1_VRSEFF_RESET = 1'h1;

// VrsConfig1.VRSO_EN
parameter VRSCONFIG1_VRSO_EN_WIDTH = 1;
parameter VRSCONFIG1_VRSO_EN_LSB = 7;
parameter VRSCONFIG1_VRSO_EN_MASK = 8'h80;
parameter VRSCONFIG1_VRSO_EN_RESET = 1'h0;


// VrsConfig2
parameter VRSCONFIG2_ADDR = 8'h2d;
parameter VRSCONFIG2_RESET = 8'h0;

// VrsConfig2.VRS_OL_DIAG
parameter VRSCONFIG2_VRS_OL_DIAG_WIDTH = 7;
parameter VRSCONFIG2_VRS_OL_DIAG_LSB = 0;
parameter VRSCONFIG2_VRS_OL_DIAG_MASK = 8'h7f;
parameter VRSCONFIG2_VRS_OL_DIAG_RESET = 7'h0;


// MscConfig0
parameter MSCCONFIG0_ADDR = 8'h2e;
parameter MSCCONFIG0_RESET = 8'h0;

// MscConfig0.MSC_CLK_DIV_CFG
parameter MSCCONFIG0_MSC_CLK_DIV_CFG_WIDTH = 3;
parameter MSCCONFIG0_MSC_CLK_DIV_CFG_LSB = 0;
parameter MSCCONFIG0_MSC_CLK_DIV_CFG_MASK = 8'h7;
parameter MSCCONFIG0_MSC_CLK_DIV_CFG_RESET = 3'h0;

// MscConfig0.MSC_SV_EN
parameter MSCCONFIG0_MSC_SV_EN_WIDTH = 1;
parameter MSCCONFIG0_MSC_SV_EN_LSB = 3;
parameter MSCCONFIG0_MSC_SV_EN_MASK = 8'h8;
parameter MSCCONFIG0_MSC_SV_EN_RESET = 1'h0;


// MscConfig1
parameter MSCCONFIG1_ADDR = 8'h2f;
parameter MSCCONFIG1_RESET = 8'h1;

// MscConfig1.MSC_CRC_CFG
parameter MSCCONFIG1_MSC_CRC_CFG_WIDTH = 1;
parameter MSCCONFIG1_MSC_CRC_CFG_LSB = 0;
parameter MSCCONFIG1_MSC_CRC_CFG_MASK = 8'h1;
parameter MSCCONFIG1_MSC_CRC_CFG_RESET = 1'h1;

// MscConfig1.MSC_UP_FRAME
parameter MSCCONFIG1_MSC_UP_FRAME_WIDTH = 1;
parameter MSCCONFIG1_MSC_UP_FRAME_LSB = 1;
parameter MSCCONFIG1_MSC_UP_FRAME_MASK = 8'h2;
parameter MSCCONFIG1_MSC_UP_FRAME_RESET = 1'h0;

// MscConfig1.MSC_ADDR_MODE
parameter MSCCONFIG1_MSC_ADDR_MODE_WIDTH = 1;
parameter MSCCONFIG1_MSC_ADDR_MODE_LSB = 2;
parameter MSCCONFIG1_MSC_ADDR_MODE_MASK = 8'h4;
parameter MSCCONFIG1_MSC_ADDR_MODE_RESET = 1'h0;

// MscConfig1.MSC_ADDR_CFG
parameter MSCCONFIG1_MSC_ADDR_CFG_WIDTH = 4;
parameter MSCCONFIG1_MSC_ADDR_CFG_LSB = 3;
parameter MSCCONFIG1_MSC_ADDR_CFG_MASK = 8'h78;
parameter MSCCONFIG1_MSC_ADDR_CFG_RESET = 4'h0;

// MscConfig1.OD_MISO
parameter MSCCONFIG1_OD_MISO_WIDTH = 1;
parameter MSCCONFIG1_OD_MISO_LSB = 7;
parameter MSCCONFIG1_OD_MISO_MASK = 8'h80;
parameter MSCCONFIG1_OD_MISO_RESET = 1'h0;


// AoutConfig
parameter AOUTCONFIG_ADDR = 8'h30;
parameter AOUTCONFIG_RESET = 8'h10;

// AoutConfig.AMUX
parameter AOUTCONFIG_AMUX_WIDTH = 4;
parameter AOUTCONFIG_AMUX_LSB = 0;
parameter AOUTCONFIG_AMUX_MASK = 8'hf;
parameter AOUTCONFIG_AMUX_RESET = 4'h0;

// AoutConfig.VDDIO_RNG
parameter AOUTCONFIG_VDDIO_RNG_WIDTH = 2;
parameter AOUTCONFIG_VDDIO_RNG_LSB = 4;
parameter AOUTCONFIG_VDDIO_RNG_MASK = 8'h30;
parameter AOUTCONFIG_VDDIO_RNG_RESET = 2'h1;

// AoutConfig.VPWR_RNG
parameter AOUTCONFIG_VPWR_RNG_WIDTH = 1;
parameter AOUTCONFIG_VPWR_RNG_LSB = 6;
parameter AOUTCONFIG_VPWR_RNG_MASK = 8'h40;
parameter AOUTCONFIG_VPWR_RNG_RESET = 1'h0;


// RstbConfig
parameter RSTBCONFIG_ADDR = 8'h31;
parameter RSTBCONFIG_RESET = 8'h7;

// RstbConfig.VDD5_UV_RSTB_CFG
parameter RSTBCONFIG_VDD5_UV_RSTB_CFG_WIDTH = 1;
parameter RSTBCONFIG_VDD5_UV_RSTB_CFG_LSB = 0;
parameter RSTBCONFIG_VDD5_UV_RSTB_CFG_MASK = 8'h1;
parameter RSTBCONFIG_VDD5_UV_RSTB_CFG_RESET = 1'h1;

// RstbConfig.VDD5_OV_RSTB_CFG
parameter RSTBCONFIG_VDD5_OV_RSTB_CFG_WIDTH = 1;
parameter RSTBCONFIG_VDD5_OV_RSTB_CFG_LSB = 1;
parameter RSTBCONFIG_VDD5_OV_RSTB_CFG_MASK = 8'h2;
parameter RSTBCONFIG_VDD5_OV_RSTB_CFG_RESET = 1'h1;

// RstbConfig.WD_RSTB_CFG
parameter RSTBCONFIG_WD_RSTB_CFG_WIDTH = 1;
parameter RSTBCONFIG_WD_RSTB_CFG_LSB = 2;
parameter RSTBCONFIG_WD_RSTB_CFG_MASK = 8'h4;
parameter RSTBCONFIG_WD_RSTB_CFG_RESET = 1'h1;


// FaultbConfig0
parameter FAULTBCONFIG0_ADDR = 8'h32;
parameter FAULTBCONFIG0_RESET = 8'h3f;

// FaultbConfig0.WD_SV_FAIL_DIAG
parameter FAULTBCONFIG0_WD_SV_FAIL_DIAG_WIDTH = 1;
parameter FAULTBCONFIG0_WD_SV_FAIL_DIAG_LSB = 0;
parameter FAULTBCONFIG0_WD_SV_FAIL_DIAG_MASK = 8'h1;
parameter FAULTBCONFIG0_WD_SV_FAIL_DIAG_RESET = 1'h1;

// FaultbConfig0.SPI_MSC_FAIL_DIAG
parameter FAULTBCONFIG0_SPI_MSC_FAIL_DIAG_WIDTH = 1;
parameter FAULTBCONFIG0_SPI_MSC_FAIL_DIAG_LSB = 1;
parameter FAULTBCONFIG0_SPI_MSC_FAIL_DIAG_MASK = 8'h2;
parameter FAULTBCONFIG0_SPI_MSC_FAIL_DIAG_RESET = 1'h1;

// FaultbConfig0.OTP_FAIL_DIAG
parameter FAULTBCONFIG0_OTP_FAIL_DIAG_WIDTH = 1;
parameter FAULTBCONFIG0_OTP_FAIL_DIAG_LSB = 2;
parameter FAULTBCONFIG0_OTP_FAIL_DIAG_MASK = 8'h4;
parameter FAULTBCONFIG0_OTP_FAIL_DIAG_RESET = 1'h1;

// FaultbConfig0.FAULT_VRS_WD_DIAG
parameter FAULTBCONFIG0_FAULT_VRS_WD_DIAG_WIDTH = 1;
parameter FAULTBCONFIG0_FAULT_VRS_WD_DIAG_LSB = 3;
parameter FAULTBCONFIG0_FAULT_VRS_WD_DIAG_MASK = 8'h8;
parameter FAULTBCONFIG0_FAULT_VRS_WD_DIAG_RESET = 1'h1;

// FaultbConfig0.VRS_OL_SC_DIAG
parameter FAULTBCONFIG0_VRS_OL_SC_DIAG_WIDTH = 1;
parameter FAULTBCONFIG0_VRS_OL_SC_DIAG_LSB = 4;
parameter FAULTBCONFIG0_VRS_OL_SC_DIAG_MASK = 8'h10;
parameter FAULTBCONFIG0_VRS_OL_SC_DIAG_RESET = 1'h1;

// FaultbConfig0.GND_FAIL_DIAG
parameter FAULTBCONFIG0_GND_FAIL_DIAG_WIDTH = 1;
parameter FAULTBCONFIG0_GND_FAIL_DIAG_LSB = 5;
parameter FAULTBCONFIG0_GND_FAIL_DIAG_MASK = 8'h20;
parameter FAULTBCONFIG0_GND_FAIL_DIAG_RESET = 1'h1;

// FaultbConfig0.FAULTB_LATCH_DATA
parameter FAULTBCONFIG0_FAULTB_LATCH_DATA_WIDTH = 1;
parameter FAULTBCONFIG0_FAULTB_LATCH_DATA_LSB = 7;
parameter FAULTBCONFIG0_FAULTB_LATCH_DATA_MASK = 8'h80;
parameter FAULTBCONFIG0_FAULTB_LATCH_DATA_RESET = 1'h0;


// FaultbConfig1
parameter FAULTBCONFIG1_ADDR = 8'h33;
parameter FAULTBCONFIG1_RESET = 8'hff;

// FaultbConfig1.SUP_REGL_DIAG
parameter FAULTBCONFIG1_SUP_REGL_DIAG_WIDTH = 1;
parameter FAULTBCONFIG1_SUP_REGL_DIAG_LSB = 0;
parameter FAULTBCONFIG1_SUP_REGL_DIAG_MASK = 8'h1;
parameter FAULTBCONFIG1_SUP_REGL_DIAG_RESET = 1'h1;

// FaultbConfig1.CP_UV_DIAG
parameter FAULTBCONFIG1_CP_UV_DIAG_WIDTH = 1;
parameter FAULTBCONFIG1_CP_UV_DIAG_LSB = 1;
parameter FAULTBCONFIG1_CP_UV_DIAG_MASK = 8'h2;
parameter FAULTBCONFIG1_CP_UV_DIAG_RESET = 1'h1;

// FaultbConfig1.VDDIO_UV_DIAG
parameter FAULTBCONFIG1_VDDIO_UV_DIAG_WIDTH = 1;
parameter FAULTBCONFIG1_VDDIO_UV_DIAG_LSB = 2;
parameter FAULTBCONFIG1_VDDIO_UV_DIAG_MASK = 8'h4;
parameter FAULTBCONFIG1_VDDIO_UV_DIAG_RESET = 1'h1;

// FaultbConfig1.VDDIO_OV_DIAG
parameter FAULTBCONFIG1_VDDIO_OV_DIAG_WIDTH = 1;
parameter FAULTBCONFIG1_VDDIO_OV_DIAG_LSB = 3;
parameter FAULTBCONFIG1_VDDIO_OV_DIAG_MASK = 8'h8;
parameter FAULTBCONFIG1_VDDIO_OV_DIAG_RESET = 1'h1;

// FaultbConfig1.VPWR_UV_DIAG
parameter FAULTBCONFIG1_VPWR_UV_DIAG_WIDTH = 1;
parameter FAULTBCONFIG1_VPWR_UV_DIAG_LSB = 4;
parameter FAULTBCONFIG1_VPWR_UV_DIAG_MASK = 8'h10;
parameter FAULTBCONFIG1_VPWR_UV_DIAG_RESET = 1'h1;

// FaultbConfig1.VPWR_OV_DIAG
parameter FAULTBCONFIG1_VPWR_OV_DIAG_WIDTH = 1;
parameter FAULTBCONFIG1_VPWR_OV_DIAG_LSB = 5;
parameter FAULTBCONFIG1_VPWR_OV_DIAG_MASK = 8'h20;
parameter FAULTBCONFIG1_VPWR_OV_DIAG_RESET = 1'h1;

// FaultbConfig1.VDD5_UV_DIAG
parameter FAULTBCONFIG1_VDD5_UV_DIAG_WIDTH = 1;
parameter FAULTBCONFIG1_VDD5_UV_DIAG_LSB = 6;
parameter FAULTBCONFIG1_VDD5_UV_DIAG_MASK = 8'h40;
parameter FAULTBCONFIG1_VDD5_UV_DIAG_RESET = 1'h1;

// FaultbConfig1.VDD5_OV_DIAG
parameter FAULTBCONFIG1_VDD5_OV_DIAG_WIDTH = 1;
parameter FAULTBCONFIG1_VDD5_OV_DIAG_LSB = 7;
parameter FAULTBCONFIG1_VDD5_OV_DIAG_MASK = 8'h80;
parameter FAULTBCONFIG1_VDD5_OV_DIAG_RESET = 1'h1;


// FaultbConfig2
parameter FAULTBCONFIG2_ADDR = 8'h34;
parameter FAULTBCONFIG2_RESET = 8'h3f;

// FaultbConfig2.OL_SC_DIAG
parameter FAULTBCONFIG2_OL_SC_DIAG_WIDTH = 1;
parameter FAULTBCONFIG2_OL_SC_DIAG_LSB = 0;
parameter FAULTBCONFIG2_OL_SC_DIAG_MASK = 8'h1;
parameter FAULTBCONFIG2_OL_SC_DIAG_RESET = 1'h1;

// FaultbConfig2.TSD_DIAG
parameter FAULTBCONFIG2_TSD_DIAG_WIDTH = 1;
parameter FAULTBCONFIG2_TSD_DIAG_LSB = 1;
parameter FAULTBCONFIG2_TSD_DIAG_MASK = 8'h2;
parameter FAULTBCONFIG2_TSD_DIAG_RESET = 1'h1;

// FaultbConfig2.OC_DIAG
parameter FAULTBCONFIG2_OC_DIAG_WIDTH = 1;
parameter FAULTBCONFIG2_OC_DIAG_LSB = 2;
parameter FAULTBCONFIG2_OC_DIAG_MASK = 8'h4;
parameter FAULTBCONFIG2_OC_DIAG_RESET = 1'h1;

// FaultbConfig2.SC_IGN_DIAG
parameter FAULTBCONFIG2_SC_IGN_DIAG_WIDTH = 1;
parameter FAULTBCONFIG2_SC_IGN_DIAG_LSB = 3;
parameter FAULTBCONFIG2_SC_IGN_DIAG_MASK = 8'h8;
parameter FAULTBCONFIG2_SC_IGN_DIAG_RESET = 1'h1;

// FaultbConfig2.OL_IGN_DIAG
parameter FAULTBCONFIG2_OL_IGN_DIAG_WIDTH = 1;
parameter FAULTBCONFIG2_OL_IGN_DIAG_LSB = 4;
parameter FAULTBCONFIG2_OL_IGN_DIAG_MASK = 8'h10;
parameter FAULTBCONFIG2_OL_IGN_DIAG_RESET = 1'h1;

// FaultbConfig2.DNDIS_DRV_DIAG
parameter FAULTBCONFIG2_DNDIS_DRV_DIAG_WIDTH = 1;
parameter FAULTBCONFIG2_DNDIS_DRV_DIAG_LSB = 5;
parameter FAULTBCONFIG2_DNDIS_DRV_DIAG_MASK = 8'h20;
parameter FAULTBCONFIG2_DNDIS_DRV_DIAG_RESET = 1'h1;

// FaultbConfig2.FAULTB_SPI_CTRL_MODE
parameter FAULTBCONFIG2_FAULTB_SPI_CTRL_MODE_WIDTH = 1;
parameter FAULTBCONFIG2_FAULTB_SPI_CTRL_MODE_LSB = 6;
parameter FAULTBCONFIG2_FAULTB_SPI_CTRL_MODE_MASK = 8'h40;
parameter FAULTBCONFIG2_FAULTB_SPI_CTRL_MODE_RESET = 1'h0;

// FaultbConfig2.FAULTB_SPI_CTRL
parameter FAULTBCONFIG2_FAULTB_SPI_CTRL_WIDTH = 1;
parameter FAULTBCONFIG2_FAULTB_SPI_CTRL_LSB = 7;
parameter FAULTBCONFIG2_FAULTB_SPI_CTRL_MASK = 8'h80;
parameter FAULTBCONFIG2_FAULTB_SPI_CTRL_RESET = 1'h0;


// VrsDiag
parameter VRSDIAG_ADDR = 8'h35;
parameter VRSDIAG_RESET = 8'h0;

// VrsDiag.FAULT_VRS_WD
parameter VRSDIAG_FAULT_VRS_WD_WIDTH = 1;
parameter VRSDIAG_FAULT_VRS_WD_LSB = 0;
parameter VRSDIAG_FAULT_VRS_WD_MASK = 8'h1;
parameter VRSDIAG_FAULT_VRS_WD_RESET = 1'h0;

// VrsDiag.VRS_SCB
parameter VRSDIAG_VRS_SCB_WIDTH = 1;
parameter VRSDIAG_VRS_SCB_LSB = 1;
parameter VRSDIAG_VRS_SCB_MASK = 8'h2;
parameter VRSDIAG_VRS_SCB_RESET = 1'h0;

// VrsDiag.VRS_SCG
parameter VRSDIAG_VRS_SCG_WIDTH = 1;
parameter VRSDIAG_VRS_SCG_LSB = 2;
parameter VRSDIAG_VRS_SCG_MASK = 8'h4;
parameter VRSDIAG_VRS_SCG_RESET = 1'h0;

// VrsDiag.VRS_OL
parameter VRSDIAG_VRS_OL_WIDTH = 1;
parameter VRSDIAG_VRS_OL_LSB = 3;
parameter VRSDIAG_VRS_OL_MASK = 8'h8;
parameter VRSDIAG_VRS_OL_RESET = 1'h0;

// VrsDiag.VRS_TH_FAULT
parameter VRSDIAG_VRS_TH_FAULT_WIDTH = 1;
parameter VRSDIAG_VRS_TH_FAULT_LSB = 4;
parameter VRSDIAG_VRS_TH_FAULT_MASK = 8'h10;
parameter VRSDIAG_VRS_TH_FAULT_RESET = 1'h0;


// SupDiag
parameter SUPDIAG_ADDR = 8'h36;
parameter SUPDIAG_RESET = 8'h0;

// SupDiag.SUP_REGL
parameter SUPDIAG_SUP_REGL_WIDTH = 1;
parameter SUPDIAG_SUP_REGL_LSB = 0;
parameter SUPDIAG_SUP_REGL_MASK = 8'h1;
parameter SUPDIAG_SUP_REGL_RESET = 1'h0;

// SupDiag.CP_UV
parameter SUPDIAG_CP_UV_WIDTH = 1;
parameter SUPDIAG_CP_UV_LSB = 1;
parameter SUPDIAG_CP_UV_MASK = 8'h2;
parameter SUPDIAG_CP_UV_RESET = 1'h0;

// SupDiag.VDDIO_UV
parameter SUPDIAG_VDDIO_UV_WIDTH = 1;
parameter SUPDIAG_VDDIO_UV_LSB = 2;
parameter SUPDIAG_VDDIO_UV_MASK = 8'h4;
parameter SUPDIAG_VDDIO_UV_RESET = 1'h0;

// SupDiag.VDDIO_OV
parameter SUPDIAG_VDDIO_OV_WIDTH = 1;
parameter SUPDIAG_VDDIO_OV_LSB = 3;
parameter SUPDIAG_VDDIO_OV_MASK = 8'h8;
parameter SUPDIAG_VDDIO_OV_RESET = 1'h0;

// SupDiag.VPWR_UV
parameter SUPDIAG_VPWR_UV_WIDTH = 1;
parameter SUPDIAG_VPWR_UV_LSB = 4;
parameter SUPDIAG_VPWR_UV_MASK = 8'h10;
parameter SUPDIAG_VPWR_UV_RESET = 1'h0;

// SupDiag.VPWR_OV
parameter SUPDIAG_VPWR_OV_WIDTH = 1;
parameter SUPDIAG_VPWR_OV_LSB = 5;
parameter SUPDIAG_VPWR_OV_MASK = 8'h20;
parameter SUPDIAG_VPWR_OV_RESET = 1'h0;

// SupDiag.VDD5_UV
parameter SUPDIAG_VDD5_UV_WIDTH = 1;
parameter SUPDIAG_VDD5_UV_LSB = 6;
parameter SUPDIAG_VDD5_UV_MASK = 8'h40;
parameter SUPDIAG_VDD5_UV_RESET = 1'h0;

// SupDiag.VDD5_OV
parameter SUPDIAG_VDD5_OV_WIDTH = 1;
parameter SUPDIAG_VDD5_OV_LSB = 7;
parameter SUPDIAG_VDD5_OV_MASK = 8'h80;
parameter SUPDIAG_VDD5_OV_RESET = 1'h0;


// ExtDiag0
parameter EXTDIAG0_ADDR = 8'h37;
parameter EXTDIAG0_RESET = 8'h0;

// ExtDiag0.MSC_SPI_ERROR
parameter EXTDIAG0_MSC_SPI_ERROR_WIDTH = 1;
parameter EXTDIAG0_MSC_SPI_ERROR_LSB = 0;
parameter EXTDIAG0_MSC_SPI_ERROR_MASK = 8'h1;
parameter EXTDIAG0_MSC_SPI_ERROR_RESET = 1'h0;

// ExtDiag0.MSC_SV_ERROR
parameter EXTDIAG0_MSC_SV_ERROR_WIDTH = 1;
parameter EXTDIAG0_MSC_SV_ERROR_LSB = 1;
parameter EXTDIAG0_MSC_SV_ERROR_MASK = 8'h2;
parameter EXTDIAG0_MSC_SV_ERROR_RESET = 1'h0;

// ExtDiag0.WD_WARN
parameter EXTDIAG0_WD_WARN_WIDTH = 1;
parameter EXTDIAG0_WD_WARN_LSB = 2;
parameter EXTDIAG0_WD_WARN_MASK = 8'h4;
parameter EXTDIAG0_WD_WARN_RESET = 1'h0;

// ExtDiag0.WD_FAIL
parameter EXTDIAG0_WD_FAIL_WIDTH = 1;
parameter EXTDIAG0_WD_FAIL_LSB = 3;
parameter EXTDIAG0_WD_FAIL_MASK = 8'h8;
parameter EXTDIAG0_WD_FAIL_RESET = 1'h0;

// ExtDiag0.FUSE_CHECK_ERROR
parameter EXTDIAG0_FUSE_CHECK_ERROR_WIDTH = 1;
parameter EXTDIAG0_FUSE_CHECK_ERROR_LSB = 4;
parameter EXTDIAG0_FUSE_CHECK_ERROR_MASK = 8'h10;
parameter EXTDIAG0_FUSE_CHECK_ERROR_RESET = 1'h0;

// ExtDiag0.OTP_USAGE_FAULT
parameter EXTDIAG0_OTP_USAGE_FAULT_WIDTH = 1;
parameter EXTDIAG0_OTP_USAGE_FAULT_LSB = 5;
parameter EXTDIAG0_OTP_USAGE_FAULT_MASK = 8'h20;
parameter EXTDIAG0_OTP_USAGE_FAULT_RESET = 1'h0;

// ExtDiag0.SELF_TEST_ERROR
parameter EXTDIAG0_SELF_TEST_ERROR_WIDTH = 1;
parameter EXTDIAG0_SELF_TEST_ERROR_LSB = 6;
parameter EXTDIAG0_SELF_TEST_ERROR_MASK = 8'h40;
parameter EXTDIAG0_SELF_TEST_ERROR_RESET = 1'h0;


// ExtDiag1
parameter EXTDIAG1_ADDR = 8'h38;
parameter EXTDIAG1_RESET = 8'h0;

// ExtDiag1.PGND_LOSS
parameter EXTDIAG1_PGND_LOSS_WIDTH = 1;
parameter EXTDIAG1_PGND_LOSS_LSB = 0;
parameter EXTDIAG1_PGND_LOSS_MASK = 8'h1;
parameter EXTDIAG1_PGND_LOSS_RESET = 1'h0;

// ExtDiag1.AGND_LOSS
parameter EXTDIAG1_AGND_LOSS_WIDTH = 1;
parameter EXTDIAG1_AGND_LOSS_LSB = 1;
parameter EXTDIAG1_AGND_LOSS_MASK = 8'h2;
parameter EXTDIAG1_AGND_LOSS_RESET = 1'h0;

// ExtDiag1.GNDIO_LOSS
parameter EXTDIAG1_GNDIO_LOSS_WIDTH = 1;
parameter EXTDIAG1_GNDIO_LOSS_LSB = 2;
parameter EXTDIAG1_GNDIO_LOSS_MASK = 8'h4;
parameter EXTDIAG1_GNDIO_LOSS_RESET = 1'h0;

// ExtDiag1.VDIG_1P5V_OV
parameter EXTDIAG1_VDIG_1P5V_OV_WIDTH = 1;
parameter EXTDIAG1_VDIG_1P5V_OV_LSB = 3;
parameter EXTDIAG1_VDIG_1P5V_OV_MASK = 8'h8;
parameter EXTDIAG1_VDIG_1P5V_OV_RESET = 1'h0;

// ExtDiag1.VDIG_1P5V_UV
parameter EXTDIAG1_VDIG_1P5V_UV_WIDTH = 1;
parameter EXTDIAG1_VDIG_1P5V_UV_LSB = 4;
parameter EXTDIAG1_VDIG_1P5V_UV_MASK = 8'h10;
parameter EXTDIAG1_VDIG_1P5V_UV_RESET = 1'h0;

// ExtDiag1.VANA_1P5V_UV
parameter EXTDIAG1_VANA_1P5V_UV_WIDTH = 1;
parameter EXTDIAG1_VANA_1P5V_UV_LSB = 5;
parameter EXTDIAG1_VANA_1P5V_UV_MASK = 8'h20;
parameter EXTDIAG1_VANA_1P5V_UV_RESET = 1'h0;

// ExtDiag1.VANA_1P5V_OV
parameter EXTDIAG1_VANA_1P5V_OV_WIDTH = 1;
parameter EXTDIAG1_VANA_1P5V_OV_LSB = 6;
parameter EXTDIAG1_VANA_1P5V_OV_MASK = 8'h40;
parameter EXTDIAG1_VANA_1P5V_OV_RESET = 1'h0;

// ExtDiag1.DIS_DRV
parameter EXTDIAG1_DIS_DRV_WIDTH = 1;
parameter EXTDIAG1_DIS_DRV_LSB = 7;
parameter EXTDIAG1_DIS_DRV_MASK = 8'h80;
parameter EXTDIAG1_DIS_DRV_RESET = 1'h0;


// InjDiag0
parameter INJDIAG0_ADDR = 8'h39;
parameter INJDIAG0_RESET = 8'h0;

// InjDiag0.SCG_INJ1
parameter INJDIAG0_SCG_INJ1_WIDTH = 1;
parameter INJDIAG0_SCG_INJ1_LSB = 0;
parameter INJDIAG0_SCG_INJ1_MASK = 8'h1;
parameter INJDIAG0_SCG_INJ1_RESET = 1'h0;

// InjDiag0.OL_INJ1
parameter INJDIAG0_OL_INJ1_WIDTH = 1;
parameter INJDIAG0_OL_INJ1_LSB = 1;
parameter INJDIAG0_OL_INJ1_MASK = 8'h2;
parameter INJDIAG0_OL_INJ1_RESET = 1'h0;

// InjDiag0.TSD_INJ1
parameter INJDIAG0_TSD_INJ1_WIDTH = 1;
parameter INJDIAG0_TSD_INJ1_LSB = 2;
parameter INJDIAG0_TSD_INJ1_MASK = 8'h4;
parameter INJDIAG0_TSD_INJ1_RESET = 1'h0;

// InjDiag0.OC_INJ1
parameter INJDIAG0_OC_INJ1_WIDTH = 1;
parameter INJDIAG0_OC_INJ1_LSB = 3;
parameter INJDIAG0_OC_INJ1_MASK = 8'h8;
parameter INJDIAG0_OC_INJ1_RESET = 1'h0;

// InjDiag0.SCG_INJ2
parameter INJDIAG0_SCG_INJ2_WIDTH = 1;
parameter INJDIAG0_SCG_INJ2_LSB = 4;
parameter INJDIAG0_SCG_INJ2_MASK = 8'h10;
parameter INJDIAG0_SCG_INJ2_RESET = 1'h0;

// InjDiag0.OL_INJ2
parameter INJDIAG0_OL_INJ2_WIDTH = 1;
parameter INJDIAG0_OL_INJ2_LSB = 5;
parameter INJDIAG0_OL_INJ2_MASK = 8'h20;
parameter INJDIAG0_OL_INJ2_RESET = 1'h0;

// InjDiag0.TSD_INJ2
parameter INJDIAG0_TSD_INJ2_WIDTH = 1;
parameter INJDIAG0_TSD_INJ2_LSB = 6;
parameter INJDIAG0_TSD_INJ2_MASK = 8'h40;
parameter INJDIAG0_TSD_INJ2_RESET = 1'h0;

// InjDiag0.OC_INJ2
parameter INJDIAG0_OC_INJ2_WIDTH = 1;
parameter INJDIAG0_OC_INJ2_LSB = 7;
parameter INJDIAG0_OC_INJ2_MASK = 8'h80;
parameter INJDIAG0_OC_INJ2_RESET = 1'h0;


// InjDiag1
parameter INJDIAG1_ADDR = 8'h3a;
parameter INJDIAG1_RESET = 8'h0;

// InjDiag1.SCG_INJ3
parameter INJDIAG1_SCG_INJ3_WIDTH = 1;
parameter INJDIAG1_SCG_INJ3_LSB = 0;
parameter INJDIAG1_SCG_INJ3_MASK = 8'h1;
parameter INJDIAG1_SCG_INJ3_RESET = 1'h0;

// InjDiag1.OL_INJ3
parameter INJDIAG1_OL_INJ3_WIDTH = 1;
parameter INJDIAG1_OL_INJ3_LSB = 1;
parameter INJDIAG1_OL_INJ3_MASK = 8'h2;
parameter INJDIAG1_OL_INJ3_RESET = 1'h0;

// InjDiag1.TSD_INJ3
parameter INJDIAG1_TSD_INJ3_WIDTH = 1;
parameter INJDIAG1_TSD_INJ3_LSB = 2;
parameter INJDIAG1_TSD_INJ3_MASK = 8'h4;
parameter INJDIAG1_TSD_INJ3_RESET = 1'h0;

// InjDiag1.OC_INJ3
parameter INJDIAG1_OC_INJ3_WIDTH = 1;
parameter INJDIAG1_OC_INJ3_LSB = 3;
parameter INJDIAG1_OC_INJ3_MASK = 8'h8;
parameter INJDIAG1_OC_INJ3_RESET = 1'h0;

// InjDiag1.SCG_INJ4
parameter INJDIAG1_SCG_INJ4_WIDTH = 1;
parameter INJDIAG1_SCG_INJ4_LSB = 4;
parameter INJDIAG1_SCG_INJ4_MASK = 8'h10;
parameter INJDIAG1_SCG_INJ4_RESET = 1'h0;

// InjDiag1.OL_INJ4
parameter INJDIAG1_OL_INJ4_WIDTH = 1;
parameter INJDIAG1_OL_INJ4_LSB = 5;
parameter INJDIAG1_OL_INJ4_MASK = 8'h20;
parameter INJDIAG1_OL_INJ4_RESET = 1'h0;

// InjDiag1.TSD_INJ4
parameter INJDIAG1_TSD_INJ4_WIDTH = 1;
parameter INJDIAG1_TSD_INJ4_LSB = 6;
parameter INJDIAG1_TSD_INJ4_MASK = 8'h40;
parameter INJDIAG1_TSD_INJ4_RESET = 1'h0;

// InjDiag1.OC_INJ4
parameter INJDIAG1_OC_INJ4_WIDTH = 1;
parameter INJDIAG1_OC_INJ4_LSB = 7;
parameter INJDIAG1_OC_INJ4_MASK = 8'h80;
parameter INJDIAG1_OC_INJ4_RESET = 1'h0;


// IgnDiag0
parameter IGNDIAG0_ADDR = 8'h3b;
parameter IGNDIAG0_RESET = 8'h0;

// IgnDiag0.SCG_IGN1
parameter IGNDIAG0_SCG_IGN1_WIDTH = 1;
parameter IGNDIAG0_SCG_IGN1_LSB = 0;
parameter IGNDIAG0_SCG_IGN1_MASK = 8'h1;
parameter IGNDIAG0_SCG_IGN1_RESET = 1'h0;

// IgnDiag0.OL_IGN1
parameter IGNDIAG0_OL_IGN1_WIDTH = 1;
parameter IGNDIAG0_OL_IGN1_LSB = 1;
parameter IGNDIAG0_OL_IGN1_MASK = 8'h2;
parameter IGNDIAG0_OL_IGN1_RESET = 1'h0;

// IgnDiag0.SCB_IGN1
parameter IGNDIAG0_SCB_IGN1_WIDTH = 1;
parameter IGNDIAG0_SCB_IGN1_LSB = 2;
parameter IGNDIAG0_SCB_IGN1_MASK = 8'h4;
parameter IGNDIAG0_SCB_IGN1_RESET = 1'h0;

// IgnDiag0.SCG_IGN2
parameter IGNDIAG0_SCG_IGN2_WIDTH = 1;
parameter IGNDIAG0_SCG_IGN2_LSB = 3;
parameter IGNDIAG0_SCG_IGN2_MASK = 8'h8;
parameter IGNDIAG0_SCG_IGN2_RESET = 1'h0;

// IgnDiag0.OL_IGN2
parameter IGNDIAG0_OL_IGN2_WIDTH = 1;
parameter IGNDIAG0_OL_IGN2_LSB = 4;
parameter IGNDIAG0_OL_IGN2_MASK = 8'h10;
parameter IGNDIAG0_OL_IGN2_RESET = 1'h0;

// IgnDiag0.SCB_IGN2
parameter IGNDIAG0_SCB_IGN2_WIDTH = 1;
parameter IGNDIAG0_SCB_IGN2_LSB = 5;
parameter IGNDIAG0_SCB_IGN2_MASK = 8'h20;
parameter IGNDIAG0_SCB_IGN2_RESET = 1'h0;

// IgnDiag0.TSD_IGN1
parameter IGNDIAG0_TSD_IGN1_WIDTH = 1;
parameter IGNDIAG0_TSD_IGN1_LSB = 6;
parameter IGNDIAG0_TSD_IGN1_MASK = 8'h40;
parameter IGNDIAG0_TSD_IGN1_RESET = 1'h0;


// IgnDiag1
parameter IGNDIAG1_ADDR = 8'h3c;
parameter IGNDIAG1_RESET = 8'h0;

// IgnDiag1.SCG_IGN3
parameter IGNDIAG1_SCG_IGN3_WIDTH = 1;
parameter IGNDIAG1_SCG_IGN3_LSB = 0;
parameter IGNDIAG1_SCG_IGN3_MASK = 8'h1;
parameter IGNDIAG1_SCG_IGN3_RESET = 1'h0;

// IgnDiag1.OL_IGN3
parameter IGNDIAG1_OL_IGN3_WIDTH = 1;
parameter IGNDIAG1_OL_IGN3_LSB = 1;
parameter IGNDIAG1_OL_IGN3_MASK = 8'h2;
parameter IGNDIAG1_OL_IGN3_RESET = 1'h0;

// IgnDiag1.SCB_IGN3
parameter IGNDIAG1_SCB_IGN3_WIDTH = 1;
parameter IGNDIAG1_SCB_IGN3_LSB = 2;
parameter IGNDIAG1_SCB_IGN3_MASK = 8'h4;
parameter IGNDIAG1_SCB_IGN3_RESET = 1'h0;

// IgnDiag1.SCG_IGN4
parameter IGNDIAG1_SCG_IGN4_WIDTH = 1;
parameter IGNDIAG1_SCG_IGN4_LSB = 3;
parameter IGNDIAG1_SCG_IGN4_MASK = 8'h8;
parameter IGNDIAG1_SCG_IGN4_RESET = 1'h0;

// IgnDiag1.OL_IGN4
parameter IGNDIAG1_OL_IGN4_WIDTH = 1;
parameter IGNDIAG1_OL_IGN4_LSB = 4;
parameter IGNDIAG1_OL_IGN4_MASK = 8'h10;
parameter IGNDIAG1_OL_IGN4_RESET = 1'h0;

// IgnDiag1.SCB_IGN4
parameter IGNDIAG1_SCB_IGN4_WIDTH = 1;
parameter IGNDIAG1_SCB_IGN4_LSB = 5;
parameter IGNDIAG1_SCB_IGN4_MASK = 8'h20;
parameter IGNDIAG1_SCB_IGN4_RESET = 1'h0;

// IgnDiag1.TSD_IGN2
parameter IGNDIAG1_TSD_IGN2_WIDTH = 1;
parameter IGNDIAG1_TSD_IGN2_LSB = 6;
parameter IGNDIAG1_TSD_IGN2_MASK = 8'h40;
parameter IGNDIAG1_TSD_IGN2_RESET = 1'h0;


// HtrDiag0
parameter HTRDIAG0_ADDR = 8'h3d;
parameter HTRDIAG0_RESET = 8'h0;

// HtrDiag0.SCG_HTR1
parameter HTRDIAG0_SCG_HTR1_WIDTH = 1;
parameter HTRDIAG0_SCG_HTR1_LSB = 0;
parameter HTRDIAG0_SCG_HTR1_MASK = 8'h1;
parameter HTRDIAG0_SCG_HTR1_RESET = 1'h0;

// HtrDiag0.OL_HTR1
parameter HTRDIAG0_OL_HTR1_WIDTH = 1;
parameter HTRDIAG0_OL_HTR1_LSB = 1;
parameter HTRDIAG0_OL_HTR1_MASK = 8'h2;
parameter HTRDIAG0_OL_HTR1_RESET = 1'h0;

// HtrDiag0.TSD_HTR1
parameter HTRDIAG0_TSD_HTR1_WIDTH = 1;
parameter HTRDIAG0_TSD_HTR1_LSB = 2;
parameter HTRDIAG0_TSD_HTR1_MASK = 8'h4;
parameter HTRDIAG0_TSD_HTR1_RESET = 1'h0;

// HtrDiag0.OC_HTR1
parameter HTRDIAG0_OC_HTR1_WIDTH = 1;
parameter HTRDIAG0_OC_HTR1_LSB = 3;
parameter HTRDIAG0_OC_HTR1_MASK = 8'h8;
parameter HTRDIAG0_OC_HTR1_RESET = 1'h0;

// HtrDiag0.SCG_HTR2
parameter HTRDIAG0_SCG_HTR2_WIDTH = 1;
parameter HTRDIAG0_SCG_HTR2_LSB = 4;
parameter HTRDIAG0_SCG_HTR2_MASK = 8'h10;
parameter HTRDIAG0_SCG_HTR2_RESET = 1'h0;

// HtrDiag0.OL_HTR2
parameter HTRDIAG0_OL_HTR2_WIDTH = 1;
parameter HTRDIAG0_OL_HTR2_LSB = 5;
parameter HTRDIAG0_OL_HTR2_MASK = 8'h20;
parameter HTRDIAG0_OL_HTR2_RESET = 1'h0;

// HtrDiag0.TSD_HTR2
parameter HTRDIAG0_TSD_HTR2_WIDTH = 1;
parameter HTRDIAG0_TSD_HTR2_LSB = 6;
parameter HTRDIAG0_TSD_HTR2_MASK = 8'h40;
parameter HTRDIAG0_TSD_HTR2_RESET = 1'h0;

// HtrDiag0.OC_HTR2
parameter HTRDIAG0_OC_HTR2_WIDTH = 1;
parameter HTRDIAG0_OC_HTR2_LSB = 7;
parameter HTRDIAG0_OC_HTR2_MASK = 8'h80;
parameter HTRDIAG0_OC_HTR2_RESET = 1'h0;


// RlyDiag0
parameter RLYDIAG0_ADDR = 8'h3e;
parameter RLYDIAG0_RESET = 8'h0;

// RlyDiag0.SCG_RLY1
parameter RLYDIAG0_SCG_RLY1_WIDTH = 1;
parameter RLYDIAG0_SCG_RLY1_LSB = 0;
parameter RLYDIAG0_SCG_RLY1_MASK = 8'h1;
parameter RLYDIAG0_SCG_RLY1_RESET = 1'h0;

// RlyDiag0.OL_RLY1
parameter RLYDIAG0_OL_RLY1_WIDTH = 1;
parameter RLYDIAG0_OL_RLY1_LSB = 1;
parameter RLYDIAG0_OL_RLY1_MASK = 8'h2;
parameter RLYDIAG0_OL_RLY1_RESET = 1'h0;

// RlyDiag0.TSD_RLY1
parameter RLYDIAG0_TSD_RLY1_WIDTH = 1;
parameter RLYDIAG0_TSD_RLY1_LSB = 2;
parameter RLYDIAG0_TSD_RLY1_MASK = 8'h4;
parameter RLYDIAG0_TSD_RLY1_RESET = 1'h0;

// RlyDiag0.OC_RLY1
parameter RLYDIAG0_OC_RLY1_WIDTH = 1;
parameter RLYDIAG0_OC_RLY1_LSB = 3;
parameter RLYDIAG0_OC_RLY1_MASK = 8'h8;
parameter RLYDIAG0_OC_RLY1_RESET = 1'h0;

// RlyDiag0.SCG_RLY2
parameter RLYDIAG0_SCG_RLY2_WIDTH = 1;
parameter RLYDIAG0_SCG_RLY2_LSB = 4;
parameter RLYDIAG0_SCG_RLY2_MASK = 8'h10;
parameter RLYDIAG0_SCG_RLY2_RESET = 1'h0;

// RlyDiag0.OL_RLY2
parameter RLYDIAG0_OL_RLY2_WIDTH = 1;
parameter RLYDIAG0_OL_RLY2_LSB = 5;
parameter RLYDIAG0_OL_RLY2_MASK = 8'h20;
parameter RLYDIAG0_OL_RLY2_RESET = 1'h0;

// RlyDiag0.TSD_RLY2
parameter RLYDIAG0_TSD_RLY2_WIDTH = 1;
parameter RLYDIAG0_TSD_RLY2_LSB = 6;
parameter RLYDIAG0_TSD_RLY2_MASK = 8'h40;
parameter RLYDIAG0_TSD_RLY2_RESET = 1'h0;

// RlyDiag0.OC_RLY2
parameter RLYDIAG0_OC_RLY2_WIDTH = 1;
parameter RLYDIAG0_OC_RLY2_LSB = 7;
parameter RLYDIAG0_OC_RLY2_MASK = 8'h80;
parameter RLYDIAG0_OC_RLY2_RESET = 1'h0;


// RlyDiag1
parameter RLYDIAG1_ADDR = 8'h3f;
parameter RLYDIAG1_RESET = 8'h0;

// RlyDiag1.SCG_RLY3
parameter RLYDIAG1_SCG_RLY3_WIDTH = 1;
parameter RLYDIAG1_SCG_RLY3_LSB = 0;
parameter RLYDIAG1_SCG_RLY3_MASK = 8'h1;
parameter RLYDIAG1_SCG_RLY3_RESET = 1'h0;

// RlyDiag1.OL_RLY3
parameter RLYDIAG1_OL_RLY3_WIDTH = 1;
parameter RLYDIAG1_OL_RLY3_LSB = 1;
parameter RLYDIAG1_OL_RLY3_MASK = 8'h2;
parameter RLYDIAG1_OL_RLY3_RESET = 1'h0;

// RlyDiag1.TSD_RLY3
parameter RLYDIAG1_TSD_RLY3_WIDTH = 1;
parameter RLYDIAG1_TSD_RLY3_LSB = 2;
parameter RLYDIAG1_TSD_RLY3_MASK = 8'h4;
parameter RLYDIAG1_TSD_RLY3_RESET = 1'h0;

// RlyDiag1.OC_RLY3
parameter RLYDIAG1_OC_RLY3_WIDTH = 1;
parameter RLYDIAG1_OC_RLY3_LSB = 3;
parameter RLYDIAG1_OC_RLY3_MASK = 8'h8;
parameter RLYDIAG1_OC_RLY3_RESET = 1'h0;

// RlyDiag1.SCG_RLY4
parameter RLYDIAG1_SCG_RLY4_WIDTH = 1;
parameter RLYDIAG1_SCG_RLY4_LSB = 4;
parameter RLYDIAG1_SCG_RLY4_MASK = 8'h10;
parameter RLYDIAG1_SCG_RLY4_RESET = 1'h0;

// RlyDiag1.OL_RLY4
parameter RLYDIAG1_OL_RLY4_WIDTH = 1;
parameter RLYDIAG1_OL_RLY4_LSB = 5;
parameter RLYDIAG1_OL_RLY4_MASK = 8'h20;
parameter RLYDIAG1_OL_RLY4_RESET = 1'h0;

// RlyDiag1.TSD_RLY4
parameter RLYDIAG1_TSD_RLY4_WIDTH = 1;
parameter RLYDIAG1_TSD_RLY4_LSB = 6;
parameter RLYDIAG1_TSD_RLY4_MASK = 8'h40;
parameter RLYDIAG1_TSD_RLY4_RESET = 1'h0;

// RlyDiag1.OC_RLY4
parameter RLYDIAG1_OC_RLY4_WIDTH = 1;
parameter RLYDIAG1_OC_RLY4_LSB = 7;
parameter RLYDIAG1_OC_RLY4_MASK = 8'h80;
parameter RLYDIAG1_OC_RLY4_RESET = 1'h0;


// RlyDiag2
parameter RLYDIAG2_ADDR = 8'h40;
parameter RLYDIAG2_RESET = 8'h0;

// RlyDiag2.SCG_RLY5
parameter RLYDIAG2_SCG_RLY5_WIDTH = 1;
parameter RLYDIAG2_SCG_RLY5_LSB = 0;
parameter RLYDIAG2_SCG_RLY5_MASK = 8'h1;
parameter RLYDIAG2_SCG_RLY5_RESET = 1'h0;

// RlyDiag2.OL_RLY5
parameter RLYDIAG2_OL_RLY5_WIDTH = 1;
parameter RLYDIAG2_OL_RLY5_LSB = 1;
parameter RLYDIAG2_OL_RLY5_MASK = 8'h2;
parameter RLYDIAG2_OL_RLY5_RESET = 1'h0;

// RlyDiag2.TSD_RLY5
parameter RLYDIAG2_TSD_RLY5_WIDTH = 1;
parameter RLYDIAG2_TSD_RLY5_LSB = 2;
parameter RLYDIAG2_TSD_RLY5_MASK = 8'h4;
parameter RLYDIAG2_TSD_RLY5_RESET = 1'h0;

// RlyDiag2.OC_RLY5
parameter RLYDIAG2_OC_RLY5_WIDTH = 1;
parameter RLYDIAG2_OC_RLY5_LSB = 3;
parameter RLYDIAG2_OC_RLY5_MASK = 8'h8;
parameter RLYDIAG2_OC_RLY5_RESET = 1'h0;

// RlyDiag2.SCG_RLY6
parameter RLYDIAG2_SCG_RLY6_WIDTH = 1;
parameter RLYDIAG2_SCG_RLY6_LSB = 4;
parameter RLYDIAG2_SCG_RLY6_MASK = 8'h10;
parameter RLYDIAG2_SCG_RLY6_RESET = 1'h0;

// RlyDiag2.OL_RLY6
parameter RLYDIAG2_OL_RLY6_WIDTH = 1;
parameter RLYDIAG2_OL_RLY6_LSB = 5;
parameter RLYDIAG2_OL_RLY6_MASK = 8'h20;
parameter RLYDIAG2_OL_RLY6_RESET = 1'h0;

// RlyDiag2.TSD_RLY6
parameter RLYDIAG2_TSD_RLY6_WIDTH = 1;
parameter RLYDIAG2_TSD_RLY6_LSB = 6;
parameter RLYDIAG2_TSD_RLY6_MASK = 8'h40;
parameter RLYDIAG2_TSD_RLY6_RESET = 1'h0;

// RlyDiag2.OC_RLY6
parameter RLYDIAG2_OC_RLY6_WIDTH = 1;
parameter RLYDIAG2_OC_RLY6_LSB = 7;
parameter RLYDIAG2_OC_RLY6_MASK = 8'h80;
parameter RLYDIAG2_OC_RLY6_RESET = 1'h0;


// RlyDiag3
parameter RLYDIAG3_ADDR = 8'h41;
parameter RLYDIAG3_RESET = 8'h0;

// RlyDiag3.SCG_RLY7
parameter RLYDIAG3_SCG_RLY7_WIDTH = 1;
parameter RLYDIAG3_SCG_RLY7_LSB = 0;
parameter RLYDIAG3_SCG_RLY7_MASK = 8'h1;
parameter RLYDIAG3_SCG_RLY7_RESET = 1'h0;

// RlyDiag3.OL_RLY7
parameter RLYDIAG3_OL_RLY7_WIDTH = 1;
parameter RLYDIAG3_OL_RLY7_LSB = 1;
parameter RLYDIAG3_OL_RLY7_MASK = 8'h2;
parameter RLYDIAG3_OL_RLY7_RESET = 1'h0;

// RlyDiag3.TSD_RLY7
parameter RLYDIAG3_TSD_RLY7_WIDTH = 1;
parameter RLYDIAG3_TSD_RLY7_LSB = 2;
parameter RLYDIAG3_TSD_RLY7_MASK = 8'h4;
parameter RLYDIAG3_TSD_RLY7_RESET = 1'h0;

// RlyDiag3.OC_RLY7
parameter RLYDIAG3_OC_RLY7_WIDTH = 1;
parameter RLYDIAG3_OC_RLY7_LSB = 3;
parameter RLYDIAG3_OC_RLY7_MASK = 8'h8;
parameter RLYDIAG3_OC_RLY7_RESET = 1'h0;

// RlyDiag3.SCG_RLY8
parameter RLYDIAG3_SCG_RLY8_WIDTH = 1;
parameter RLYDIAG3_SCG_RLY8_LSB = 4;
parameter RLYDIAG3_SCG_RLY8_MASK = 8'h10;
parameter RLYDIAG3_SCG_RLY8_RESET = 1'h0;

// RlyDiag3.OL_RLY8
parameter RLYDIAG3_OL_RLY8_WIDTH = 1;
parameter RLYDIAG3_OL_RLY8_LSB = 5;
parameter RLYDIAG3_OL_RLY8_MASK = 8'h20;
parameter RLYDIAG3_OL_RLY8_RESET = 1'h0;

// RlyDiag3.TSD_RLY8
parameter RLYDIAG3_TSD_RLY8_WIDTH = 1;
parameter RLYDIAG3_TSD_RLY8_LSB = 6;
parameter RLYDIAG3_TSD_RLY8_MASK = 8'h40;
parameter RLYDIAG3_TSD_RLY8_RESET = 1'h0;

// RlyDiag3.OC_RLY8
parameter RLYDIAG3_OC_RLY8_WIDTH = 1;
parameter RLYDIAG3_OC_RLY8_LSB = 7;
parameter RLYDIAG3_OC_RLY8_MASK = 8'h80;
parameter RLYDIAG3_OC_RLY8_RESET = 1'h0;


// RlyDiag4
parameter RLYDIAG4_ADDR = 8'h42;
parameter RLYDIAG4_RESET = 8'h0;

// RlyDiag4.SCG_RLY9
parameter RLYDIAG4_SCG_RLY9_WIDTH = 1;
parameter RLYDIAG4_SCG_RLY9_LSB = 0;
parameter RLYDIAG4_SCG_RLY9_MASK = 8'h1;
parameter RLYDIAG4_SCG_RLY9_RESET = 1'h0;

// RlyDiag4.OL_RLY9
parameter RLYDIAG4_OL_RLY9_WIDTH = 1;
parameter RLYDIAG4_OL_RLY9_LSB = 1;
parameter RLYDIAG4_OL_RLY9_MASK = 8'h2;
parameter RLYDIAG4_OL_RLY9_RESET = 1'h0;

// RlyDiag4.TSD_RLY9
parameter RLYDIAG4_TSD_RLY9_WIDTH = 1;
parameter RLYDIAG4_TSD_RLY9_LSB = 2;
parameter RLYDIAG4_TSD_RLY9_MASK = 8'h4;
parameter RLYDIAG4_TSD_RLY9_RESET = 1'h0;

// RlyDiag4.OC_RLY9
parameter RLYDIAG4_OC_RLY9_WIDTH = 1;
parameter RLYDIAG4_OC_RLY9_LSB = 3;
parameter RLYDIAG4_OC_RLY9_MASK = 8'h8;
parameter RLYDIAG4_OC_RLY9_RESET = 1'h0;

// RlyDiag4.SCG_VLV1
parameter RLYDIAG4_SCG_VLV1_WIDTH = 1;
parameter RLYDIAG4_SCG_VLV1_LSB = 4;
parameter RLYDIAG4_SCG_VLV1_MASK = 8'h10;
parameter RLYDIAG4_SCG_VLV1_RESET = 1'h0;

// RlyDiag4.OL_VLV1
parameter RLYDIAG4_OL_VLV1_WIDTH = 1;
parameter RLYDIAG4_OL_VLV1_LSB = 5;
parameter RLYDIAG4_OL_VLV1_MASK = 8'h20;
parameter RLYDIAG4_OL_VLV1_RESET = 1'h0;

// RlyDiag4.TSD_VLV1
parameter RLYDIAG4_TSD_VLV1_WIDTH = 1;
parameter RLYDIAG4_TSD_VLV1_LSB = 6;
parameter RLYDIAG4_TSD_VLV1_MASK = 8'h40;
parameter RLYDIAG4_TSD_VLV1_RESET = 1'h0;

// RlyDiag4.OC_VLV1
parameter RLYDIAG4_OC_VLV1_WIDTH = 1;
parameter RLYDIAG4_OC_VLV1_LSB = 7;
parameter RLYDIAG4_OC_VLV1_MASK = 8'h80;
parameter RLYDIAG4_OC_VLV1_RESET = 1'h0;


// VlvDiag
parameter VLVDIAG_ADDR = 8'h43;
parameter VLVDIAG_RESET = 8'h0;

// VlvDiag.SCG_VLV2
parameter VLVDIAG_SCG_VLV2_WIDTH = 1;
parameter VLVDIAG_SCG_VLV2_LSB = 0;
parameter VLVDIAG_SCG_VLV2_MASK = 8'h1;
parameter VLVDIAG_SCG_VLV2_RESET = 1'h0;

// VlvDiag.OL_VLV2
parameter VLVDIAG_OL_VLV2_WIDTH = 1;
parameter VLVDIAG_OL_VLV2_LSB = 1;
parameter VLVDIAG_OL_VLV2_MASK = 8'h2;
parameter VLVDIAG_OL_VLV2_RESET = 1'h0;

// VlvDiag.TSD_VLV2
parameter VLVDIAG_TSD_VLV2_WIDTH = 1;
parameter VLVDIAG_TSD_VLV2_LSB = 2;
parameter VLVDIAG_TSD_VLV2_MASK = 8'h4;
parameter VLVDIAG_TSD_VLV2_RESET = 1'h0;

// VlvDiag.OC_VLV2
parameter VLVDIAG_OC_VLV2_WIDTH = 1;
parameter VLVDIAG_OC_VLV2_LSB = 3;
parameter VLVDIAG_OC_VLV2_MASK = 8'h8;
parameter VLVDIAG_OC_VLV2_RESET = 1'h0;

// VlvDiag.SCG_VLV3
parameter VLVDIAG_SCG_VLV3_WIDTH = 1;
parameter VLVDIAG_SCG_VLV3_LSB = 4;
parameter VLVDIAG_SCG_VLV3_MASK = 8'h10;
parameter VLVDIAG_SCG_VLV3_RESET = 1'h0;

// VlvDiag.OL_VLV3
parameter VLVDIAG_OL_VLV3_WIDTH = 1;
parameter VLVDIAG_OL_VLV3_LSB = 5;
parameter VLVDIAG_OL_VLV3_MASK = 8'h20;
parameter VLVDIAG_OL_VLV3_RESET = 1'h0;

// VlvDiag.TSD_VLV3
parameter VLVDIAG_TSD_VLV3_WIDTH = 1;
parameter VLVDIAG_TSD_VLV3_LSB = 6;
parameter VLVDIAG_TSD_VLV3_MASK = 8'h40;
parameter VLVDIAG_TSD_VLV3_RESET = 1'h0;

// VlvDiag.OC_VLV3
parameter VLVDIAG_OC_VLV3_WIDTH = 1;
parameter VLVDIAG_OC_VLV3_LSB = 7;
parameter VLVDIAG_OC_VLV3_MASK = 8'h80;
parameter VLVDIAG_OC_VLV3_RESET = 1'h0;


// HbDiag0
parameter HBDIAG0_ADDR = 8'h44;
parameter HBDIAG0_RESET = 8'h0;

// HbDiag0.TSD_HS1
parameter HBDIAG0_TSD_HS1_WIDTH = 1;
parameter HBDIAG0_TSD_HS1_LSB = 0;
parameter HBDIAG0_TSD_HS1_MASK = 8'h1;
parameter HBDIAG0_TSD_HS1_RESET = 1'h0;

// HbDiag0.OC_HS1
parameter HBDIAG0_OC_HS1_WIDTH = 1;
parameter HBDIAG0_OC_HS1_LSB = 1;
parameter HBDIAG0_OC_HS1_MASK = 8'h2;
parameter HBDIAG0_OC_HS1_RESET = 1'h0;

// HbDiag0.TSD_LS1
parameter HBDIAG0_TSD_LS1_WIDTH = 1;
parameter HBDIAG0_TSD_LS1_LSB = 2;
parameter HBDIAG0_TSD_LS1_MASK = 8'h4;
parameter HBDIAG0_TSD_LS1_RESET = 1'h0;

// HbDiag0.OC_LS1
parameter HBDIAG0_OC_LS1_WIDTH = 1;
parameter HBDIAG0_OC_LS1_LSB = 3;
parameter HBDIAG0_OC_LS1_MASK = 8'h8;
parameter HBDIAG0_OC_LS1_RESET = 1'h0;

// HbDiag0.SCG_HB1
parameter HBDIAG0_SCG_HB1_WIDTH = 1;
parameter HBDIAG0_SCG_HB1_LSB = 4;
parameter HBDIAG0_SCG_HB1_MASK = 8'h10;
parameter HBDIAG0_SCG_HB1_RESET = 1'h0;

// HbDiag0.SCB_HB1
parameter HBDIAG0_SCB_HB1_WIDTH = 1;
parameter HBDIAG0_SCB_HB1_LSB = 5;
parameter HBDIAG0_SCB_HB1_MASK = 8'h20;
parameter HBDIAG0_SCB_HB1_RESET = 1'h0;

// HbDiag0.OL_HB1
parameter HBDIAG0_OL_HB1_WIDTH = 1;
parameter HBDIAG0_OL_HB1_LSB = 6;
parameter HBDIAG0_OL_HB1_MASK = 8'h40;
parameter HBDIAG0_OL_HB1_RESET = 1'h0;


// HbDiag1
parameter HBDIAG1_ADDR = 8'h45;
parameter HBDIAG1_RESET = 8'h0;

// HbDiag1.TSD_HS2
parameter HBDIAG1_TSD_HS2_WIDTH = 1;
parameter HBDIAG1_TSD_HS2_LSB = 0;
parameter HBDIAG1_TSD_HS2_MASK = 8'h1;
parameter HBDIAG1_TSD_HS2_RESET = 1'h0;

// HbDiag1.OC_HS2
parameter HBDIAG1_OC_HS2_WIDTH = 1;
parameter HBDIAG1_OC_HS2_LSB = 1;
parameter HBDIAG1_OC_HS2_MASK = 8'h2;
parameter HBDIAG1_OC_HS2_RESET = 1'h0;

// HbDiag1.TSD_LS2
parameter HBDIAG1_TSD_LS2_WIDTH = 1;
parameter HBDIAG1_TSD_LS2_LSB = 2;
parameter HBDIAG1_TSD_LS2_MASK = 8'h4;
parameter HBDIAG1_TSD_LS2_RESET = 1'h0;

// HbDiag1.OC_LS2
parameter HBDIAG1_OC_LS2_WIDTH = 1;
parameter HBDIAG1_OC_LS2_LSB = 3;
parameter HBDIAG1_OC_LS2_MASK = 8'h8;
parameter HBDIAG1_OC_LS2_RESET = 1'h0;

// HbDiag1.SCG_HB2
parameter HBDIAG1_SCG_HB2_WIDTH = 1;
parameter HBDIAG1_SCG_HB2_LSB = 4;
parameter HBDIAG1_SCG_HB2_MASK = 8'h10;
parameter HBDIAG1_SCG_HB2_RESET = 1'h0;

// HbDiag1.SCB_HB2
parameter HBDIAG1_SCB_HB2_WIDTH = 1;
parameter HBDIAG1_SCB_HB2_LSB = 5;
parameter HBDIAG1_SCB_HB2_MASK = 8'h20;
parameter HBDIAG1_SCB_HB2_RESET = 1'h0;

// HbDiag1.OL_HB2
parameter HBDIAG1_OL_HB2_WIDTH = 1;
parameter HBDIAG1_OL_HB2_LSB = 6;
parameter HBDIAG1_OL_HB2_MASK = 8'h40;
parameter HBDIAG1_OL_HB2_RESET = 1'h0;


// RstDiag
parameter RSTDIAG_ADDR = 8'h46;
parameter RSTDIAG_RESET = 8'h0;

// RstDiag.RSTB_EVENT
parameter RSTDIAG_RSTB_EVENT_WIDTH = 1;
parameter RSTDIAG_RSTB_EVENT_LSB = 0;
parameter RSTDIAG_RSTB_EVENT_MASK = 8'h1;
parameter RSTDIAG_RSTB_EVENT_RESET = 1'h0;

// RstDiag.WD_RST_EVENT
parameter RSTDIAG_WD_RST_EVENT_WIDTH = 1;
parameter RSTDIAG_WD_RST_EVENT_LSB = 1;
parameter RSTDIAG_WD_RST_EVENT_MASK = 8'h2;
parameter RSTDIAG_WD_RST_EVENT_RESET = 1'h0;

// RstDiag.SOFTWARE_RST_EVENT
parameter RSTDIAG_SOFTWARE_RST_EVENT_WIDTH = 1;
parameter RSTDIAG_SOFTWARE_RST_EVENT_LSB = 2;
parameter RSTDIAG_SOFTWARE_RST_EVENT_MASK = 8'h4;
parameter RSTDIAG_SOFTWARE_RST_EVENT_RESET = 1'h0;

// RstDiag.VDD5_UV_RST_EVENT
parameter RSTDIAG_VDD5_UV_RST_EVENT_WIDTH = 1;
parameter RSTDIAG_VDD5_UV_RST_EVENT_LSB = 3;
parameter RSTDIAG_VDD5_UV_RST_EVENT_MASK = 8'h8;
parameter RSTDIAG_VDD5_UV_RST_EVENT_RESET = 1'h0;

// RstDiag.VDD5_OV_RST_EVENT
parameter RSTDIAG_VDD5_OV_RST_EVENT_WIDTH = 1;
parameter RSTDIAG_VDD5_OV_RST_EVENT_LSB = 4;
parameter RSTDIAG_VDD5_OV_RST_EVENT_MASK = 8'h10;
parameter RSTDIAG_VDD5_OV_RST_EVENT_RESET = 1'h0;

// RstDiag.POR_EVENT
parameter RSTDIAG_POR_EVENT_WIDTH = 1;
parameter RSTDIAG_POR_EVENT_LSB = 5;
parameter RSTDIAG_POR_EVENT_MASK = 8'h20;
parameter RSTDIAG_POR_EVENT_RESET = 1'h0;


// GLBStatus
parameter GLBSTATUS_ADDR = 8'h47;
parameter GLBSTATUS_RESET = 8'h0;

// GLBStatus.TSD_OC_FAIL
parameter GLBSTATUS_TSD_OC_FAIL_WIDTH = 1;
parameter GLBSTATUS_TSD_OC_FAIL_LSB = 0;
parameter GLBSTATUS_TSD_OC_FAIL_MASK = 8'h1;
parameter GLBSTATUS_TSD_OC_FAIL_RESET = 1'h0;

// GLBStatus.SC_OL_FAIL
parameter GLBSTATUS_SC_OL_FAIL_WIDTH = 1;
parameter GLBSTATUS_SC_OL_FAIL_LSB = 1;
parameter GLBSTATUS_SC_OL_FAIL_MASK = 8'h2;
parameter GLBSTATUS_SC_OL_FAIL_RESET = 1'h0;

// GLBStatus.WD_SV_FAIL
parameter GLBSTATUS_WD_SV_FAIL_WIDTH = 1;
parameter GLBSTATUS_WD_SV_FAIL_LSB = 2;
parameter GLBSTATUS_WD_SV_FAIL_MASK = 8'h4;
parameter GLBSTATUS_WD_SV_FAIL_RESET = 1'h0;

// GLBStatus.SUP_FAIL_DIS_DRV
parameter GLBSTATUS_SUP_FAIL_DIS_DRV_WIDTH = 1;
parameter GLBSTATUS_SUP_FAIL_DIS_DRV_LSB = 3;
parameter GLBSTATUS_SUP_FAIL_DIS_DRV_MASK = 8'h8;
parameter GLBSTATUS_SUP_FAIL_DIS_DRV_RESET = 1'h0;

// GLBStatus.VRS_FAIL
parameter GLBSTATUS_VRS_FAIL_WIDTH = 1;
parameter GLBSTATUS_VRS_FAIL_LSB = 4;
parameter GLBSTATUS_VRS_FAIL_MASK = 8'h10;
parameter GLBSTATUS_VRS_FAIL_RESET = 1'h0;

// GLBStatus.OTP_FAIL
parameter GLBSTATUS_OTP_FAIL_WIDTH = 1;
parameter GLBSTATUS_OTP_FAIL_LSB = 5;
parameter GLBSTATUS_OTP_FAIL_MASK = 8'h20;
parameter GLBSTATUS_OTP_FAIL_RESET = 1'h0;

// GLBStatus.SPI_MSC_FAIL
parameter GLBSTATUS_SPI_MSC_FAIL_WIDTH = 1;
parameter GLBSTATUS_SPI_MSC_FAIL_LSB = 6;
parameter GLBSTATUS_SPI_MSC_FAIL_MASK = 8'h40;
parameter GLBSTATUS_SPI_MSC_FAIL_RESET = 1'h0;

// GLBStatus.GND_FAIL
parameter GLBSTATUS_GND_FAIL_WIDTH = 1;
parameter GLBSTATUS_GND_FAIL_LSB = 7;
parameter GLBSTATUS_GND_FAIL_MASK = 8'h80;
parameter GLBSTATUS_GND_FAIL_RESET = 1'h0;


// WdQuestion
parameter WDQUESTION_ADDR = 8'h48;
parameter WDQUESTION_RESET = 8'h0;

// WdQuestion.LFSR
parameter WDQUESTION_LFSR_WIDTH = 8;
parameter WDQUESTION_LFSR_LSB = 0;
parameter WDQUESTION_LFSR_MASK = 8'hff;
parameter WDQUESTION_LFSR_RESET = 8'h0;


// WdPassCnt
parameter WDPASSCNT_ADDR = 8'h49;
parameter WDPASSCNT_RESET = 8'h0;

// WdPassCnt.WD_RFH_CNT
parameter WDPASSCNT_WD_RFH_CNT_WIDTH = 3;
parameter WDPASSCNT_WD_RFH_CNT_LSB = 0;
parameter WDPASSCNT_WD_RFH_CNT_MASK = 8'h7;
parameter WDPASSCNT_WD_RFH_CNT_RESET = 3'h0;


// WdFailCnt
parameter WDFAILCNT_ADDR = 8'h4a;
parameter WDFAILCNT_RESET = 8'h0;

// WdFailCnt.WD_ERR_CNT
parameter WDFAILCNT_WD_ERR_CNT_WIDTH = 3;
parameter WDFAILCNT_WD_ERR_CNT_LSB = 0;
parameter WDFAILCNT_WD_ERR_CNT_MASK = 8'h7;
parameter WDFAILCNT_WD_ERR_CNT_RESET = 3'h0;

// WdFailCnt.RST_ERR_CNT
parameter WDFAILCNT_RST_ERR_CNT_WIDTH = 3;
parameter WDFAILCNT_RST_ERR_CNT_LSB = 3;
parameter WDFAILCNT_RST_ERR_CNT_MASK = 8'h38;
parameter WDFAILCNT_RST_ERR_CNT_RESET = 3'h0;


// PSState0
parameter PSSTATE0_ADDR = 8'h4b;
parameter PSSTATE0_RESET = 8'h0;

// PSState0.OUT_STATE_IGN
parameter PSSTATE0_OUT_STATE_IGN_WIDTH = 4;
parameter PSSTATE0_OUT_STATE_IGN_LSB = 0;
parameter PSSTATE0_OUT_STATE_IGN_MASK = 8'hf;
parameter PSSTATE0_OUT_STATE_IGN_RESET = 4'h0;

// PSState0.OUT_STATE_INJ
parameter PSSTATE0_OUT_STATE_INJ_WIDTH = 4;
parameter PSSTATE0_OUT_STATE_INJ_LSB = 4;
parameter PSSTATE0_OUT_STATE_INJ_MASK = 8'hf0;
parameter PSSTATE0_OUT_STATE_INJ_RESET = 4'h0;


// PSState1
parameter PSSTATE1_ADDR = 8'h4c;
parameter PSSTATE1_RESET = 8'h0;

// PSState1.OUT_STATE_RLY
parameter PSSTATE1_OUT_STATE_RLY_WIDTH = 8;
parameter PSSTATE1_OUT_STATE_RLY_LSB = 0;
parameter PSSTATE1_OUT_STATE_RLY_MASK = 8'hff;
parameter PSSTATE1_OUT_STATE_RLY_RESET = 8'h0;


// PSState2
parameter PSSTATE2_ADDR = 8'h4d;
parameter PSSTATE2_RESET = 8'h0;

// PSState2.OUT_STATE_RLY
parameter PSSTATE2_OUT_STATE_RLY_WIDTH = 1;
parameter PSSTATE2_OUT_STATE_RLY_LSB = 0;
parameter PSSTATE2_OUT_STATE_RLY_MASK = 8'h1;
parameter PSSTATE2_OUT_STATE_RLY_RESET = 1'h0;

// PSState2.OUT_STATE_HTR
parameter PSSTATE2_OUT_STATE_HTR_WIDTH = 2;
parameter PSSTATE2_OUT_STATE_HTR_LSB = 1;
parameter PSSTATE2_OUT_STATE_HTR_MASK = 8'h6;
parameter PSSTATE2_OUT_STATE_HTR_RESET = 2'h0;

// PSState2.OUT_STATE_VLV
parameter PSSTATE2_OUT_STATE_VLV_WIDTH = 3;
parameter PSSTATE2_OUT_STATE_VLV_LSB = 3;
parameter PSSTATE2_OUT_STATE_VLV_MASK = 8'h38;
parameter PSSTATE2_OUT_STATE_VLV_RESET = 3'h0;


// PSState3
parameter PSSTATE3_ADDR = 8'h4e;
parameter PSSTATE3_RESET = 8'h0;

// PSState3.OUT_STATE_HS
parameter PSSTATE3_OUT_STATE_HS_WIDTH = 2;
parameter PSSTATE3_OUT_STATE_HS_LSB = 0;
parameter PSSTATE3_OUT_STATE_HS_MASK = 8'h3;
parameter PSSTATE3_OUT_STATE_HS_RESET = 2'h0;

// PSState3.OUT_STATE_LS
parameter PSSTATE3_OUT_STATE_LS_WIDTH = 2;
parameter PSSTATE3_OUT_STATE_LS_LSB = 2;
parameter PSSTATE3_OUT_STATE_LS_MASK = 8'hc;
parameter PSSTATE3_OUT_STATE_LS_RESET = 2'h0;


// InState0
parameter INSTATE0_ADDR = 8'h4f;
parameter INSTATE0_RESET = 8'h0;

// InState0.DIN
parameter INSTATE0_DIN_WIDTH = 8;
parameter INSTATE0_DIN_LSB = 0;
parameter INSTATE0_DIN_MASK = 8'hff;
parameter INSTATE0_DIN_RESET = 8'h0;


// InState1
parameter INSTATE1_ADDR = 8'h50;
parameter INSTATE1_RESET = 8'h0;

// InState1.DIN
parameter INSTATE1_DIN_WIDTH = 5;
parameter INSTATE1_DIN_LSB = 0;
parameter INSTATE1_DIN_MASK = 8'h1f;
parameter INSTATE1_DIN_RESET = 5'h0;


// EnState0
parameter ENSTATE0_ADDR = 8'h51;
parameter ENSTATE0_RESET = 8'h0;

// EnState0.OE
parameter ENSTATE0_OE_WIDTH = 1;
parameter ENSTATE0_OE_LSB = 0;
parameter ENSTATE0_OE_MASK = 8'h1;
parameter ENSTATE0_OE_RESET = 1'h0;

// EnState0.DEN_RLY
parameter ENSTATE0_DEN_RLY_WIDTH = 1;
parameter ENSTATE0_DEN_RLY_LSB = 1;
parameter ENSTATE0_DEN_RLY_MASK = 8'h2;
parameter ENSTATE0_DEN_RLY_RESET = 1'h0;

// EnState0.DEN_DRV
parameter ENSTATE0_DEN_DRV_WIDTH = 1;
parameter ENSTATE0_DEN_DRV_LSB = 2;
parameter ENSTATE0_DEN_DRV_MASK = 8'h4;
parameter ENSTATE0_DEN_DRV_RESET = 1'h0;

// EnState0.DNDIS_DRV
parameter ENSTATE0_DNDIS_DRV_WIDTH = 1;
parameter ENSTATE0_DNDIS_DRV_LSB = 3;
parameter ENSTATE0_DNDIS_DRV_MASK = 8'h8;
parameter ENSTATE0_DNDIS_DRV_RESET = 1'h0;


// MaskID
parameter MASKID_ADDR = 8'h52;
parameter MASKID_RESET = 8'h0;

// MaskID.MASK_ID
parameter MASKID_MASK_ID_WIDTH = 5;
parameter MASKID_MASK_ID_LSB = 0;
parameter MASKID_MASK_ID_MASK = 8'h1f;
parameter MASKID_MASK_ID_RESET = 5'h0;


// Cmd0
parameter CMD0_ADDR = 8'h53;
parameter CMD0_RESET = 8'h0;

// Cmd0.Code
parameter CMD0_CODE_WIDTH = 8;
parameter CMD0_CODE_LSB = 0;
parameter CMD0_CODE_MASK = 8'hff;
parameter CMD0_CODE_RESET = 8'h0;


// CmdWdCheck
parameter CMDWDCHECK_ADDR = 8'h54;
parameter CMDWDCHECK_RESET = 8'h0;

// CmdWdCheck.MCU_REPLY
parameter CMDWDCHECK_MCU_REPLY_WIDTH = 8;
parameter CMDWDCHECK_MCU_REPLY_LSB = 0;
parameter CMDWDCHECK_MCU_REPLY_MASK = 8'hff;
parameter CMDWDCHECK_MCU_REPLY_RESET = 8'h0;


// CmdWdLdSd
parameter CMDWDLDSD_ADDR = 8'h55;
parameter CMDWDLDSD_RESET = 8'h0;

// CmdWdLdSd.SEED
parameter CMDWDLDSD_SEED_WIDTH = 8;
parameter CMDWDLDSD_SEED_LSB = 0;
parameter CMDWDLDSD_SEED_MASK = 8'hff;
parameter CMDWDLDSD_SEED_RESET = 8'h0;


// CmdSoftRst
parameter CMDSOFTRST_ADDR = 8'h56;
parameter CMDSOFTRST_RESET = 8'h0;

// CmdSoftRst.SOFTWARE_RST
parameter CMDSOFTRST_SOFTWARE_RST_WIDTH = 8;
parameter CMDSOFTRST_SOFTWARE_RST_LSB = 0;
parameter CMDSOFTRST_SOFTWARE_RST_MASK = 8'hff;
parameter CMDSOFTRST_SOFTWARE_RST_RESET = 8'h0;


// MscRCmd0
parameter MSCRCMD0_ADDR = 8'h57;
parameter MSCRCMD0_RESET = 8'h0;

// MscRCmd0.DisDrvConfig0
parameter MSCRCMD0_DISDRVCONFIG0_WIDTH = 1;
parameter MSCRCMD0_DISDRVCONFIG0_LSB = 0;
parameter MSCRCMD0_DISDRVCONFIG0_MASK = 8'h1;
parameter MSCRCMD0_DISDRVCONFIG0_RESET = 1'h0;

// MscRCmd0.DisDrvConfig1
parameter MSCRCMD0_DISDRVCONFIG1_WIDTH = 1;
parameter MSCRCMD0_DISDRVCONFIG1_LSB = 1;
parameter MSCRCMD0_DISDRVCONFIG1_MASK = 8'h2;
parameter MSCRCMD0_DISDRVCONFIG1_RESET = 1'h0;

// MscRCmd0.DisDrvConfig2
parameter MSCRCMD0_DISDRVCONFIG2_WIDTH = 1;
parameter MSCRCMD0_DISDRVCONFIG2_LSB = 2;
parameter MSCRCMD0_DISDRVCONFIG2_MASK = 8'h4;
parameter MSCRCMD0_DISDRVCONFIG2_RESET = 1'h0;

// MscRCmd0.DenConfig0
parameter MSCRCMD0_DENCONFIG0_WIDTH = 1;
parameter MSCRCMD0_DENCONFIG0_LSB = 3;
parameter MSCRCMD0_DENCONFIG0_MASK = 8'h8;
parameter MSCRCMD0_DENCONFIG0_RESET = 1'h0;

// MscRCmd0.DenConfig1
parameter MSCRCMD0_DENCONFIG1_WIDTH = 1;
parameter MSCRCMD0_DENCONFIG1_LSB = 4;
parameter MSCRCMD0_DENCONFIG1_MASK = 8'h10;
parameter MSCRCMD0_DENCONFIG1_RESET = 1'h0;

// MscRCmd0.DenConfig2
parameter MSCRCMD0_DENCONFIG2_WIDTH = 1;
parameter MSCRCMD0_DENCONFIG2_LSB = 5;
parameter MSCRCMD0_DENCONFIG2_MASK = 8'h20;
parameter MSCRCMD0_DENCONFIG2_RESET = 1'h0;

// MscRCmd0.DenConfig3
parameter MSCRCMD0_DENCONFIG3_WIDTH = 1;
parameter MSCRCMD0_DENCONFIG3_LSB = 6;
parameter MSCRCMD0_DENCONFIG3_MASK = 8'h40;
parameter MSCRCMD0_DENCONFIG3_RESET = 1'h0;

// MscRCmd0.DenConfig4
parameter MSCRCMD0_DENCONFIG4_WIDTH = 1;
parameter MSCRCMD0_DENCONFIG4_LSB = 7;
parameter MSCRCMD0_DENCONFIG4_MASK = 8'h80;
parameter MSCRCMD0_DENCONFIG4_RESET = 1'h0;


// MscRCmd1
parameter MSCRCMD1_ADDR = 8'h58;
parameter MSCRCMD1_RESET = 8'h0;

// MscRCmd1.OEConfig0
parameter MSCRCMD1_OECONFIG0_WIDTH = 1;
parameter MSCRCMD1_OECONFIG0_LSB = 0;
parameter MSCRCMD1_OECONFIG0_MASK = 8'h1;
parameter MSCRCMD1_OECONFIG0_RESET = 1'h0;

// MscRCmd1.OEConfig1
parameter MSCRCMD1_OECONFIG1_WIDTH = 1;
parameter MSCRCMD1_OECONFIG1_LSB = 1;
parameter MSCRCMD1_OECONFIG1_MASK = 8'h2;
parameter MSCRCMD1_OECONFIG1_RESET = 1'h0;

// MscRCmd1.OEConfig2
parameter MSCRCMD1_OECONFIG2_WIDTH = 1;
parameter MSCRCMD1_OECONFIG2_LSB = 2;
parameter MSCRCMD1_OECONFIG2_MASK = 8'h4;
parameter MSCRCMD1_OECONFIG2_RESET = 1'h0;

// MscRCmd1.OEConfig3
parameter MSCRCMD1_OECONFIG3_WIDTH = 1;
parameter MSCRCMD1_OECONFIG3_LSB = 3;
parameter MSCRCMD1_OECONFIG3_MASK = 8'h8;
parameter MSCRCMD1_OECONFIG3_RESET = 1'h0;

// MscRCmd1.Cont0
parameter MSCRCMD1_CONT0_WIDTH = 1;
parameter MSCRCMD1_CONT0_LSB = 4;
parameter MSCRCMD1_CONT0_MASK = 8'h10;
parameter MSCRCMD1_CONT0_RESET = 1'h0;

// MscRCmd1.Cont1
parameter MSCRCMD1_CONT1_WIDTH = 1;
parameter MSCRCMD1_CONT1_LSB = 5;
parameter MSCRCMD1_CONT1_MASK = 8'h20;
parameter MSCRCMD1_CONT1_RESET = 1'h0;

// MscRCmd1.Cont2
parameter MSCRCMD1_CONT2_WIDTH = 1;
parameter MSCRCMD1_CONT2_LSB = 6;
parameter MSCRCMD1_CONT2_MASK = 8'h40;
parameter MSCRCMD1_CONT2_RESET = 1'h0;


// MscRCmd2
parameter MSCRCMD2_ADDR = 8'h59;
parameter MSCRCMD2_RESET = 8'h0;

// MscRCmd2.DDConfig0
parameter MSCRCMD2_DDCONFIG0_WIDTH = 1;
parameter MSCRCMD2_DDCONFIG0_LSB = 0;
parameter MSCRCMD2_DDCONFIG0_MASK = 8'h1;
parameter MSCRCMD2_DDCONFIG0_RESET = 1'h0;

// MscRCmd2.DDConfig1
parameter MSCRCMD2_DDCONFIG1_WIDTH = 1;
parameter MSCRCMD2_DDCONFIG1_LSB = 1;
parameter MSCRCMD2_DDCONFIG1_MASK = 8'h2;
parameter MSCRCMD2_DDCONFIG1_RESET = 1'h0;

// MscRCmd2.DDConfig2
parameter MSCRCMD2_DDCONFIG2_WIDTH = 1;
parameter MSCRCMD2_DDCONFIG2_LSB = 2;
parameter MSCRCMD2_DDCONFIG2_MASK = 8'h4;
parameter MSCRCMD2_DDCONFIG2_RESET = 1'h0;

// MscRCmd2.BRIConfig
parameter MSCRCMD2_BRICONFIG_WIDTH = 1;
parameter MSCRCMD2_BRICONFIG_LSB = 3;
parameter MSCRCMD2_BRICONFIG_MASK = 8'h8;
parameter MSCRCMD2_BRICONFIG_RESET = 1'h0;

// MscRCmd2.DlyOffConfig
parameter MSCRCMD2_DLYOFFCONFIG_WIDTH = 1;
parameter MSCRCMD2_DLYOFFCONFIG_LSB = 4;
parameter MSCRCMD2_DLYOFFCONFIG_MASK = 8'h10;
parameter MSCRCMD2_DLYOFFCONFIG_RESET = 1'h0;

// MscRCmd2.CurrLimConfig0
parameter MSCRCMD2_CURRLIMCONFIG0_WIDTH = 1;
parameter MSCRCMD2_CURRLIMCONFIG0_LSB = 5;
parameter MSCRCMD2_CURRLIMCONFIG0_MASK = 8'h20;
parameter MSCRCMD2_CURRLIMCONFIG0_RESET = 1'h0;

// MscRCmd2.CurrLimConfig1
parameter MSCRCMD2_CURRLIMCONFIG1_WIDTH = 1;
parameter MSCRCMD2_CURRLIMCONFIG1_LSB = 6;
parameter MSCRCMD2_CURRLIMCONFIG1_MASK = 8'h40;
parameter MSCRCMD2_CURRLIMCONFIG1_RESET = 1'h0;

// MscRCmd2.CurrLimConfig2
parameter MSCRCMD2_CURRLIMCONFIG2_WIDTH = 1;
parameter MSCRCMD2_CURRLIMCONFIG2_LSB = 7;
parameter MSCRCMD2_CURRLIMCONFIG2_MASK = 8'h80;
parameter MSCRCMD2_CURRLIMCONFIG2_RESET = 1'h0;


// MscRCmd3
parameter MSCRCMD3_ADDR = 8'h5a;
parameter MSCRCMD3_RESET = 8'h0;

// MscRCmd3.OutDiagConfig0
parameter MSCRCMD3_OUTDIAGCONFIG0_WIDTH = 1;
parameter MSCRCMD3_OUTDIAGCONFIG0_LSB = 0;
parameter MSCRCMD3_OUTDIAGCONFIG0_MASK = 8'h1;
parameter MSCRCMD3_OUTDIAGCONFIG0_RESET = 1'h0;

// MscRCmd3.OutDiagConfig1
parameter MSCRCMD3_OUTDIAGCONFIG1_WIDTH = 1;
parameter MSCRCMD3_OUTDIAGCONFIG1_LSB = 1;
parameter MSCRCMD3_OUTDIAGCONFIG1_MASK = 8'h2;
parameter MSCRCMD3_OUTDIAGCONFIG1_RESET = 1'h0;

// MscRCmd3.OutDiagConfig2
parameter MSCRCMD3_OUTDIAGCONFIG2_WIDTH = 1;
parameter MSCRCMD3_OUTDIAGCONFIG2_LSB = 2;
parameter MSCRCMD3_OUTDIAGCONFIG2_MASK = 8'h4;
parameter MSCRCMD3_OUTDIAGCONFIG2_RESET = 1'h0;

// MscRCmd3.OutDiagConfig3
parameter MSCRCMD3_OUTDIAGCONFIG3_WIDTH = 1;
parameter MSCRCMD3_OUTDIAGCONFIG3_LSB = 3;
parameter MSCRCMD3_OUTDIAGCONFIG3_MASK = 8'h8;
parameter MSCRCMD3_OUTDIAGCONFIG3_RESET = 1'h0;

// MscRCmd3.OutDiagConfig4
parameter MSCRCMD3_OUTDIAGCONFIG4_WIDTH = 1;
parameter MSCRCMD3_OUTDIAGCONFIG4_LSB = 4;
parameter MSCRCMD3_OUTDIAGCONFIG4_MASK = 8'h10;
parameter MSCRCMD3_OUTDIAGCONFIG4_RESET = 1'h0;

// MscRCmd3.IgnDiagConfig
parameter MSCRCMD3_IGNDIAGCONFIG_WIDTH = 1;
parameter MSCRCMD3_IGNDIAGCONFIG_LSB = 5;
parameter MSCRCMD3_IGNDIAGCONFIG_MASK = 8'h20;
parameter MSCRCMD3_IGNDIAGCONFIG_RESET = 1'h0;


// MscRCmd4
parameter MSCRCMD4_ADDR = 8'h5b;
parameter MSCRCMD4_RESET = 8'h0;

// MscRCmd4.DinConfig0
parameter MSCRCMD4_DINCONFIG0_WIDTH = 1;
parameter MSCRCMD4_DINCONFIG0_LSB = 0;
parameter MSCRCMD4_DINCONFIG0_MASK = 8'h1;
parameter MSCRCMD4_DINCONFIG0_RESET = 1'h0;

// MscRCmd4.DinConfig1
parameter MSCRCMD4_DINCONFIG1_WIDTH = 1;
parameter MSCRCMD4_DINCONFIG1_LSB = 1;
parameter MSCRCMD4_DINCONFIG1_MASK = 8'h2;
parameter MSCRCMD4_DINCONFIG1_RESET = 1'h0;

// MscRCmd4.DinConfig2
parameter MSCRCMD4_DINCONFIG2_WIDTH = 1;
parameter MSCRCMD4_DINCONFIG2_LSB = 2;
parameter MSCRCMD4_DINCONFIG2_MASK = 8'h4;
parameter MSCRCMD4_DINCONFIG2_RESET = 1'h0;

// MscRCmd4.DinConfig3
parameter MSCRCMD4_DINCONFIG3_WIDTH = 1;
parameter MSCRCMD4_DINCONFIG3_LSB = 3;
parameter MSCRCMD4_DINCONFIG3_MASK = 8'h8;
parameter MSCRCMD4_DINCONFIG3_RESET = 1'h0;

// MscRCmd4.DinConfig4
parameter MSCRCMD4_DINCONFIG4_WIDTH = 1;
parameter MSCRCMD4_DINCONFIG4_LSB = 4;
parameter MSCRCMD4_DINCONFIG4_MASK = 8'h10;
parameter MSCRCMD4_DINCONFIG4_RESET = 1'h0;

// MscRCmd4.DinConfig5
parameter MSCRCMD4_DINCONFIG5_WIDTH = 1;
parameter MSCRCMD4_DINCONFIG5_LSB = 5;
parameter MSCRCMD4_DINCONFIG5_MASK = 8'h20;
parameter MSCRCMD4_DINCONFIG5_RESET = 1'h0;

// MscRCmd4.DinConfig6
parameter MSCRCMD4_DINCONFIG6_WIDTH = 1;
parameter MSCRCMD4_DINCONFIG6_LSB = 6;
parameter MSCRCMD4_DINCONFIG6_MASK = 8'h40;
parameter MSCRCMD4_DINCONFIG6_RESET = 1'h0;

// MscRCmd4.DinConfig7
parameter MSCRCMD4_DINCONFIG7_WIDTH = 1;
parameter MSCRCMD4_DINCONFIG7_LSB = 7;
parameter MSCRCMD4_DINCONFIG7_MASK = 8'h80;
parameter MSCRCMD4_DINCONFIG7_RESET = 1'h0;


// MscRCmd5
parameter MSCRCMD5_ADDR = 8'h5c;
parameter MSCRCMD5_RESET = 8'h0;

// MscRCmd5.DinConfig8
parameter MSCRCMD5_DINCONFIG8_WIDTH = 1;
parameter MSCRCMD5_DINCONFIG8_LSB = 0;
parameter MSCRCMD5_DINCONFIG8_MASK = 8'h1;
parameter MSCRCMD5_DINCONFIG8_RESET = 1'h0;

// MscRCmd5.DinConfig9
parameter MSCRCMD5_DINCONFIG9_WIDTH = 1;
parameter MSCRCMD5_DINCONFIG9_LSB = 1;
parameter MSCRCMD5_DINCONFIG9_MASK = 8'h2;
parameter MSCRCMD5_DINCONFIG9_RESET = 1'h0;

// MscRCmd5.DinConfig10
parameter MSCRCMD5_DINCONFIG10_WIDTH = 1;
parameter MSCRCMD5_DINCONFIG10_LSB = 2;
parameter MSCRCMD5_DINCONFIG10_MASK = 8'h4;
parameter MSCRCMD5_DINCONFIG10_RESET = 1'h0;

// MscRCmd5.DinConfig11
parameter MSCRCMD5_DINCONFIG11_WIDTH = 1;
parameter MSCRCMD5_DINCONFIG11_LSB = 3;
parameter MSCRCMD5_DINCONFIG11_MASK = 8'h8;
parameter MSCRCMD5_DINCONFIG11_RESET = 1'h0;

// MscRCmd5.RstbConfig
parameter MSCRCMD5_RSTBCONFIG_WIDTH = 1;
parameter MSCRCMD5_RSTBCONFIG_LSB = 4;
parameter MSCRCMD5_RSTBCONFIG_MASK = 8'h10;
parameter MSCRCMD5_RSTBCONFIG_RESET = 1'h0;

// MscRCmd5.FaultbConfig0
parameter MSCRCMD5_FAULTBCONFIG0_WIDTH = 1;
parameter MSCRCMD5_FAULTBCONFIG0_LSB = 5;
parameter MSCRCMD5_FAULTBCONFIG0_MASK = 8'h20;
parameter MSCRCMD5_FAULTBCONFIG0_RESET = 1'h0;

// MscRCmd5.FaultbConfig1
parameter MSCRCMD5_FAULTBCONFIG1_WIDTH = 1;
parameter MSCRCMD5_FAULTBCONFIG1_LSB = 6;
parameter MSCRCMD5_FAULTBCONFIG1_MASK = 8'h40;
parameter MSCRCMD5_FAULTBCONFIG1_RESET = 1'h0;

// MscRCmd5.FaultbConfig2
parameter MSCRCMD5_FAULTBCONFIG2_WIDTH = 1;
parameter MSCRCMD5_FAULTBCONFIG2_LSB = 7;
parameter MSCRCMD5_FAULTBCONFIG2_MASK = 8'h80;
parameter MSCRCMD5_FAULTBCONFIG2_RESET = 1'h0;


// MscRCmd6
parameter MSCRCMD6_ADDR = 8'h5d;
parameter MSCRCMD6_RESET = 8'h0;

// MscRCmd6.WDConfig0
parameter MSCRCMD6_WDCONFIG0_WIDTH = 1;
parameter MSCRCMD6_WDCONFIG0_LSB = 0;
parameter MSCRCMD6_WDCONFIG0_MASK = 8'h1;
parameter MSCRCMD6_WDCONFIG0_RESET = 1'h0;

// MscRCmd6.WDConfig1
parameter MSCRCMD6_WDCONFIG1_WIDTH = 1;
parameter MSCRCMD6_WDCONFIG1_LSB = 1;
parameter MSCRCMD6_WDCONFIG1_MASK = 8'h2;
parameter MSCRCMD6_WDCONFIG1_RESET = 1'h0;

// MscRCmd6.VrsConfig0
parameter MSCRCMD6_VRSCONFIG0_WIDTH = 1;
parameter MSCRCMD6_VRSCONFIG0_LSB = 2;
parameter MSCRCMD6_VRSCONFIG0_MASK = 8'h4;
parameter MSCRCMD6_VRSCONFIG0_RESET = 1'h0;

// MscRCmd6.VrsConfig1
parameter MSCRCMD6_VRSCONFIG1_WIDTH = 1;
parameter MSCRCMD6_VRSCONFIG1_LSB = 3;
parameter MSCRCMD6_VRSCONFIG1_MASK = 8'h8;
parameter MSCRCMD6_VRSCONFIG1_RESET = 1'h0;

// MscRCmd6.VrsConfig2
parameter MSCRCMD6_VRSCONFIG2_WIDTH = 1;
parameter MSCRCMD6_VRSCONFIG2_LSB = 4;
parameter MSCRCMD6_VRSCONFIG2_MASK = 8'h10;
parameter MSCRCMD6_VRSCONFIG2_RESET = 1'h0;

// MscRCmd6.MscConfig0
parameter MSCRCMD6_MSCCONFIG0_WIDTH = 1;
parameter MSCRCMD6_MSCCONFIG0_LSB = 5;
parameter MSCRCMD6_MSCCONFIG0_MASK = 8'h20;
parameter MSCRCMD6_MSCCONFIG0_RESET = 1'h0;

// MscRCmd6.MscConfig1
parameter MSCRCMD6_MSCCONFIG1_WIDTH = 1;
parameter MSCRCMD6_MSCCONFIG1_LSB = 6;
parameter MSCRCMD6_MSCCONFIG1_MASK = 8'h40;
parameter MSCRCMD6_MSCCONFIG1_RESET = 1'h0;

// MscRCmd6.AoutConfig
parameter MSCRCMD6_AOUTCONFIG_WIDTH = 1;
parameter MSCRCMD6_AOUTCONFIG_LSB = 7;
parameter MSCRCMD6_AOUTCONFIG_MASK = 8'h80;
parameter MSCRCMD6_AOUTCONFIG_RESET = 1'h0;


// MscRCmd7
parameter MSCRCMD7_ADDR = 8'h5e;
parameter MSCRCMD7_RESET = 8'h0;

// MscRCmd7.VrsDiag
parameter MSCRCMD7_VRSDIAG_WIDTH = 1;
parameter MSCRCMD7_VRSDIAG_LSB = 0;
parameter MSCRCMD7_VRSDIAG_MASK = 8'h1;
parameter MSCRCMD7_VRSDIAG_RESET = 1'h0;

// MscRCmd7.SupDiag
parameter MSCRCMD7_SUPDIAG_WIDTH = 1;
parameter MSCRCMD7_SUPDIAG_LSB = 1;
parameter MSCRCMD7_SUPDIAG_MASK = 8'h2;
parameter MSCRCMD7_SUPDIAG_RESET = 1'h0;

// MscRCmd7.ExtDiag0
parameter MSCRCMD7_EXTDIAG0_WIDTH = 1;
parameter MSCRCMD7_EXTDIAG0_LSB = 2;
parameter MSCRCMD7_EXTDIAG0_MASK = 8'h4;
parameter MSCRCMD7_EXTDIAG0_RESET = 1'h0;

// MscRCmd7.ExtDiag1
parameter MSCRCMD7_EXTDIAG1_WIDTH = 1;
parameter MSCRCMD7_EXTDIAG1_LSB = 3;
parameter MSCRCMD7_EXTDIAG1_MASK = 8'h8;
parameter MSCRCMD7_EXTDIAG1_RESET = 1'h0;


// MscRCmd8
parameter MSCRCMD8_ADDR = 8'h5f;
parameter MSCRCMD8_RESET = 8'h0;

// MscRCmd8.InjDiag0
parameter MSCRCMD8_INJDIAG0_WIDTH = 1;
parameter MSCRCMD8_INJDIAG0_LSB = 0;
parameter MSCRCMD8_INJDIAG0_MASK = 8'h1;
parameter MSCRCMD8_INJDIAG0_RESET = 1'h0;

// MscRCmd8.InjDiag1
parameter MSCRCMD8_INJDIAG1_WIDTH = 1;
parameter MSCRCMD8_INJDIAG1_LSB = 1;
parameter MSCRCMD8_INJDIAG1_MASK = 8'h2;
parameter MSCRCMD8_INJDIAG1_RESET = 1'h0;

// MscRCmd8.IgnDiag0
parameter MSCRCMD8_IGNDIAG0_WIDTH = 1;
parameter MSCRCMD8_IGNDIAG0_LSB = 2;
parameter MSCRCMD8_IGNDIAG0_MASK = 8'h4;
parameter MSCRCMD8_IGNDIAG0_RESET = 1'h0;

// MscRCmd8.IgnDiag1
parameter MSCRCMD8_IGNDIAG1_WIDTH = 1;
parameter MSCRCMD8_IGNDIAG1_LSB = 3;
parameter MSCRCMD8_IGNDIAG1_MASK = 8'h8;
parameter MSCRCMD8_IGNDIAG1_RESET = 1'h0;

// MscRCmd8.HbDiag0
parameter MSCRCMD8_HBDIAG0_WIDTH = 1;
parameter MSCRCMD8_HBDIAG0_LSB = 4;
parameter MSCRCMD8_HBDIAG0_MASK = 8'h10;
parameter MSCRCMD8_HBDIAG0_RESET = 1'h0;

// MscRCmd8.HbDiag1
parameter MSCRCMD8_HBDIAG1_WIDTH = 1;
parameter MSCRCMD8_HBDIAG1_LSB = 5;
parameter MSCRCMD8_HBDIAG1_MASK = 8'h20;
parameter MSCRCMD8_HBDIAG1_RESET = 1'h0;


// MscRCmd9
parameter MSCRCMD9_ADDR = 8'h60;
parameter MSCRCMD9_RESET = 8'h0;

// MscRCmd9.RlyDiag0
parameter MSCRCMD9_RLYDIAG0_WIDTH = 1;
parameter MSCRCMD9_RLYDIAG0_LSB = 0;
parameter MSCRCMD9_RLYDIAG0_MASK = 8'h1;
parameter MSCRCMD9_RLYDIAG0_RESET = 1'h0;

// MscRCmd9.RlyDiag1
parameter MSCRCMD9_RLYDIAG1_WIDTH = 1;
parameter MSCRCMD9_RLYDIAG1_LSB = 1;
parameter MSCRCMD9_RLYDIAG1_MASK = 8'h2;
parameter MSCRCMD9_RLYDIAG1_RESET = 1'h0;

// MscRCmd9.RlyDiag2
parameter MSCRCMD9_RLYDIAG2_WIDTH = 1;
parameter MSCRCMD9_RLYDIAG2_LSB = 2;
parameter MSCRCMD9_RLYDIAG2_MASK = 8'h4;
parameter MSCRCMD9_RLYDIAG2_RESET = 1'h0;

// MscRCmd9.RlyDiag3
parameter MSCRCMD9_RLYDIAG3_WIDTH = 1;
parameter MSCRCMD9_RLYDIAG3_LSB = 3;
parameter MSCRCMD9_RLYDIAG3_MASK = 8'h8;
parameter MSCRCMD9_RLYDIAG3_RESET = 1'h0;

// MscRCmd9.RlyDiag4
parameter MSCRCMD9_RLYDIAG4_WIDTH = 1;
parameter MSCRCMD9_RLYDIAG4_LSB = 4;
parameter MSCRCMD9_RLYDIAG4_MASK = 8'h10;
parameter MSCRCMD9_RLYDIAG4_RESET = 1'h0;

// MscRCmd9.HtrDiag0
parameter MSCRCMD9_HTRDIAG0_WIDTH = 1;
parameter MSCRCMD9_HTRDIAG0_LSB = 5;
parameter MSCRCMD9_HTRDIAG0_MASK = 8'h20;
parameter MSCRCMD9_HTRDIAG0_RESET = 1'h0;

// MscRCmd9.VlvDiag
parameter MSCRCMD9_VLVDIAG_WIDTH = 1;
parameter MSCRCMD9_VLVDIAG_LSB = 6;
parameter MSCRCMD9_VLVDIAG_MASK = 8'h40;
parameter MSCRCMD9_VLVDIAG_RESET = 1'h0;

// MscRCmd9.RstDiag
parameter MSCRCMD9_RSTDIAG_WIDTH = 1;
parameter MSCRCMD9_RSTDIAG_LSB = 7;
parameter MSCRCMD9_RSTDIAG_MASK = 8'h80;
parameter MSCRCMD9_RSTDIAG_RESET = 1'h0;


// MscRCmd10
parameter MSCRCMD10_ADDR = 8'h61;
parameter MSCRCMD10_RESET = 8'h0;

// MscRCmd10.GLBStatus
parameter MSCRCMD10_GLBSTATUS_WIDTH = 1;
parameter MSCRCMD10_GLBSTATUS_LSB = 0;
parameter MSCRCMD10_GLBSTATUS_MASK = 8'h1;
parameter MSCRCMD10_GLBSTATUS_RESET = 1'h0;

// MscRCmd10.WdQuestion
parameter MSCRCMD10_WDQUESTION_WIDTH = 1;
parameter MSCRCMD10_WDQUESTION_LSB = 1;
parameter MSCRCMD10_WDQUESTION_MASK = 8'h2;
parameter MSCRCMD10_WDQUESTION_RESET = 1'h0;

// MscRCmd10.WdPassCnt
parameter MSCRCMD10_WDPASSCNT_WIDTH = 1;
parameter MSCRCMD10_WDPASSCNT_LSB = 2;
parameter MSCRCMD10_WDPASSCNT_MASK = 8'h4;
parameter MSCRCMD10_WDPASSCNT_RESET = 1'h0;

// MscRCmd10.WdFailCnt
parameter MSCRCMD10_WDFAILCNT_WIDTH = 1;
parameter MSCRCMD10_WDFAILCNT_LSB = 3;
parameter MSCRCMD10_WDFAILCNT_MASK = 8'h8;
parameter MSCRCMD10_WDFAILCNT_RESET = 1'h0;


// MscRCmd11
parameter MSCRCMD11_ADDR = 8'h62;
parameter MSCRCMD11_RESET = 8'h0;

// MscRCmd11.PSState0
parameter MSCRCMD11_PSSTATE0_WIDTH = 1;
parameter MSCRCMD11_PSSTATE0_LSB = 0;
parameter MSCRCMD11_PSSTATE0_MASK = 8'h1;
parameter MSCRCMD11_PSSTATE0_RESET = 1'h0;

// MscRCmd11.PSState1
parameter MSCRCMD11_PSSTATE1_WIDTH = 1;
parameter MSCRCMD11_PSSTATE1_LSB = 1;
parameter MSCRCMD11_PSSTATE1_MASK = 8'h2;
parameter MSCRCMD11_PSSTATE1_RESET = 1'h0;

// MscRCmd11.PSState2
parameter MSCRCMD11_PSSTATE2_WIDTH = 1;
parameter MSCRCMD11_PSSTATE2_LSB = 2;
parameter MSCRCMD11_PSSTATE2_MASK = 8'h4;
parameter MSCRCMD11_PSSTATE2_RESET = 1'h0;

// MscRCmd11.PSState3
parameter MSCRCMD11_PSSTATE3_WIDTH = 1;
parameter MSCRCMD11_PSSTATE3_LSB = 3;
parameter MSCRCMD11_PSSTATE3_MASK = 8'h8;
parameter MSCRCMD11_PSSTATE3_RESET = 1'h0;

// MscRCmd11.InState0
parameter MSCRCMD11_INSTATE0_WIDTH = 1;
parameter MSCRCMD11_INSTATE0_LSB = 4;
parameter MSCRCMD11_INSTATE0_MASK = 8'h10;
parameter MSCRCMD11_INSTATE0_RESET = 1'h0;

// MscRCmd11.InState1
parameter MSCRCMD11_INSTATE1_WIDTH = 1;
parameter MSCRCMD11_INSTATE1_LSB = 5;
parameter MSCRCMD11_INSTATE1_MASK = 8'h20;
parameter MSCRCMD11_INSTATE1_RESET = 1'h0;

// MscRCmd11.EnState0
parameter MSCRCMD11_ENSTATE0_WIDTH = 1;
parameter MSCRCMD11_ENSTATE0_LSB = 6;
parameter MSCRCMD11_ENSTATE0_MASK = 8'h40;
parameter MSCRCMD11_ENSTATE0_RESET = 1'h0;

// MscRCmd11.MaskId
parameter MSCRCMD11_MASKID_WIDTH = 1;
parameter MSCRCMD11_MASKID_LSB = 7;
parameter MSCRCMD11_MASKID_MASK = 8'h80;
parameter MSCRCMD11_MASKID_RESET = 1'h0;


// CmdSpecialMode
parameter CMDSPECIALMODE_ADDR = 8'h7d;
parameter CMDSPECIALMODE_RESET = 8'h0;

// CmdSpecialMode.SM_DIS_TSD
parameter CMDSPECIALMODE_SM_DIS_TSD_WIDTH = 1;
parameter CMDSPECIALMODE_SM_DIS_TSD_LSB = 0;
parameter CMDSPECIALMODE_SM_DIS_TSD_MASK = 8'h1;
parameter CMDSPECIALMODE_SM_DIS_TSD_RESET = 1'h0;

// CmdSpecialMode.SM_DIS_VDD5_UV
parameter CMDSPECIALMODE_SM_DIS_VDD5_UV_WIDTH = 1;
parameter CMDSPECIALMODE_SM_DIS_VDD5_UV_LSB = 1;
parameter CMDSPECIALMODE_SM_DIS_VDD5_UV_MASK = 8'h2;
parameter CMDSPECIALMODE_SM_DIS_VDD5_UV_RESET = 1'h0;

// CmdSpecialMode.SM_DIS_VDD5_OV
parameter CMDSPECIALMODE_SM_DIS_VDD5_OV_WIDTH = 1;
parameter CMDSPECIALMODE_SM_DIS_VDD5_OV_LSB = 2;
parameter CMDSPECIALMODE_SM_DIS_VDD5_OV_MASK = 8'h4;
parameter CMDSPECIALMODE_SM_DIS_VDD5_OV_RESET = 1'h0;

// CmdSpecialMode.SM_DIS_VPWR_OV
parameter CMDSPECIALMODE_SM_DIS_VPWR_OV_WIDTH = 1;
parameter CMDSPECIALMODE_SM_DIS_VPWR_OV_LSB = 3;
parameter CMDSPECIALMODE_SM_DIS_VPWR_OV_MASK = 8'h8;
parameter CMDSPECIALMODE_SM_DIS_VPWR_OV_RESET = 1'h0;

// CmdSpecialMode.SM_DIS_VPWR_UV
parameter CMDSPECIALMODE_SM_DIS_VPWR_UV_WIDTH = 1;
parameter CMDSPECIALMODE_SM_DIS_VPWR_UV_LSB = 4;
parameter CMDSPECIALMODE_SM_DIS_VPWR_UV_MASK = 8'h10;
parameter CMDSPECIALMODE_SM_DIS_VPWR_UV_RESET = 1'h0;

// CmdSpecialMode.SM_DIS_VCP_UV
parameter CMDSPECIALMODE_SM_DIS_VCP_UV_WIDTH = 1;
parameter CMDSPECIALMODE_SM_DIS_VCP_UV_LSB = 5;
parameter CMDSPECIALMODE_SM_DIS_VCP_UV_MASK = 8'h20;
parameter CMDSPECIALMODE_SM_DIS_VCP_UV_RESET = 1'h0;

// CmdSpecialMode.SM_DIS_OC
parameter CMDSPECIALMODE_SM_DIS_OC_WIDTH = 1;
parameter CMDSPECIALMODE_SM_DIS_OC_LSB = 6;
parameter CMDSPECIALMODE_SM_DIS_OC_MASK = 8'h40;
parameter CMDSPECIALMODE_SM_DIS_OC_RESET = 1'h0;

// CmdSpecialMode.SM_DIS_IGN_SCG_GNDLOSS
parameter CMDSPECIALMODE_SM_DIS_IGN_SCG_GNDLOSS_WIDTH = 1;
parameter CMDSPECIALMODE_SM_DIS_IGN_SCG_GNDLOSS_LSB = 7;
parameter CMDSPECIALMODE_SM_DIS_IGN_SCG_GNDLOSS_MASK = 8'h80;
parameter CMDSPECIALMODE_SM_DIS_IGN_SCG_GNDLOSS_RESET = 1'h0;


// CmdTM
parameter CMDTM_ADDR = 8'h7e;
parameter CMDTM_RESET = 8'h0;

// CmdTM.TM_CODE
parameter CMDTM_TM_CODE_WIDTH = 8;
parameter CMDTM_TM_CODE_LSB = 0;
parameter CMDTM_TM_CODE_MASK = 8'hff;
parameter CMDTM_TM_CODE_RESET = 8'h0;


// PageVrb
parameter PAGEVRB_ADDR = 8'h7f;
parameter PAGEVRB_RESET = 8'h0;

// PageVrb.CODE
parameter PAGEVRB_CODE_WIDTH = 8;
parameter PAGEVRB_CODE_LSB = 0;
parameter PAGEVRB_CODE_MASK = 8'hff;
parameter PAGEVRB_CODE_RESET = 8'h0;


endpackage